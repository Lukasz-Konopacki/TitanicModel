���     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�	estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.3.0�ub�n_estimators�K�estimator_params�(hhhhhhhhhht��base_estimator��
deprecated��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�sqrt�hNhG        hG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h+�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�Pclass��Sex��Age��SibSp��Parch��Fare��Embarked�et�b�n_features_in_�K�
n_outputs_�K�classes_�h*h-K ��h/��R�(KK��h4�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�
estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh&hNhJ�
hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h4�f8�����R�(KhMNNNJ����J����K t�b�C              �?�t�bhQh(�scalar���hLC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hK�
node_count�M�nodes�h*h-K ��h/��R�(KM��h4�V64�����R�(Kh8N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples��missing_go_to_left�t�}�(h}hLK ��h~hLK��hhLK��h�h]K��h�h]K ��h�hLK(��h�h]K0��h�h4�u1�����R�(Kh8NNNJ����J����K t�bK8��uK@KKt�b�B@E         �                     @"��p�?�           8�@     �Y@       u                    �?.y0��k�?�            �s@���         "                    �?Hث3���?�            @m@ 4��                             �?     ��?)             P@4��                          0�FF@�'N��?&            �N@ W��                           s�,@�q�����?             9@ ���  ������������������������       �                     @�4��         	                 �܅3@8�A�0��?             6@ W��  ������������������������       �                     @        
                        p�i@@�\��N��?             3@                                  �?��
ц��?	             *@                                   �?      �?             @        ������������������������       �                     �?                                  �H@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @                                  �<@և���X�?             @ �  ������������������������       �                     @PT��  ������������������������       �                     @�U��                             �?�q�q�?             @Z��  ������������������������       �                     @0\��  ������������������������       �                      @@^��                             �?�����H�?             B@P��  ������������������������       �                     9@����                          p"�X@���|���?             &@���                            �8@؇���X�?             @ ���  ������������������������       �                     �?����  ������������������������       �                     @ ���                             �?      �?             @ ���  ������������������������       �                     �? ���  ������������������������       �                     @����          !                    �?�q�q�?             @���  ������������������������       �                      @      @������������������������       �                     �?      @#       &                   �9@���Q��?i            @e@        $       %                    �?��s����?             5@      @������������������������       �                     @        ������������������������       �                     1@        '       f                  x#J@p�B<F]�?[            �b@     @(       G                     �?��c`��?L            �^@        )       >                   �>@8����?              G@     @*       +                    �?��
ц��?             :@       @������������������������       �                     @        ,       -                   �<@�q�q�?             5@       @������������������������       �                     @       @.       =                    R@�<ݚ�?             2@    �A@/       0                 03:@@�0�!��?             1@      :@������������������������       �                     @       @1       <                   �J@���!pc�?	             &@       2       3                 03k:@      �?              @      "@������������������������       �                     �?       @4       ;                    H@����X�?             @       5       :                 X��B@r�q��?             @     @6       7                 `fF<@      �?             @      &@������������������������       �                      @       @8       9                 �|Y=@      �?              @        ������������������������       �                     �?       @������������������������       �                     �?        ������������������������       �                      @      @������������������������       �                     �?      @������������������������       �                     @      �?������������������������       �                     �?        ?       @                 `f~I@ףp=
�?             4@     @������������������������       �                     (@      @A       B                 `��I@      �?              @        ������������������������       �                     �?       C       D                 03�I@؇���X�?             @        ������������������������       �                     �?        E       F                    �?r�q��?             @        ������������������������       �                     �?       ������������������������       �                     @        H       e                    >@&:~�Q�?,             S@       I       X                    �?�Y�R_�?+            �Q@        J       K                   @B@ �o_��?             9@        ������������������������       �                     "@        L       S                    -@     ��?             0@       M       P                   �'@      �?              @        N       O                   �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        Q       R                    D@�q�q�?             @        ������������������������       �                     @       ������������������������       �                      @        T       W                   �H@      �?              @       U       V                   �E@      �?             @        ������������������������       �                      @       ������������������������       �                      @       ������������������������       �                     @        Y       d                    �?���}<S�?             G@       Z       c                   @A@��-�=��?            �C@        [       b                   �@@������?
             1@       \       ]                 �|Y=@�r����?	             .@        ������������������������       �                     @        ^       _                   �'@�<ݚ�?             "@       ������������������������       �                     @        `       a                 �|�=@�q�q�?             @        ������������������������       �                      @       ������������������������       �                     �?        ������������������������       �                      @       ������������������������       �                     6@        ������������������������       �                     @       ������������������������       �                     @        g       t                 03�U@PN��T'�?             ;@       h       i                    <@��s����?             5@        ������������������������       �                     @        j       k                    ?@      �?	             0@        ������������������������       �                     �?        l       m                    B@z�G�z�?             .@        ������������������������       �                     @        n       o                    C@�z�G��?             $@        ������������������������       �                      @        p       q                    �?      �?              @        ������������������������       �                     @       r       s                 0� Q@      �?             @        ������������������������       �                     @        ������������������������       �                     �?       ������������������������       �                     @       v       w                    :@���B���?3            �S@        ������������������������       �        
             1@       x                          �8@�jTM��?)            �N@        y       ~                    @�g�y��?             ?@        z       {                 ��W@      �?             @        ������������������������       �                      @        |       }                 �(\�?      �?              @        ������������������������       �                     �?       ������������������������       �                     �?       ������������������������       �                     ;@       �       �                    �?��S���?             >@       �       �                  DT@�ՙ/�?             5@       �       �                     �?�n_Y�K�?	             *@ ���  �       �                 X�,D@      �?             @ ���  ������������������������       �                     �?�z��  ������������������������       �                     @    t   �       �                    �?X�<ݚ�?             "@    )   ������������������������       �                     @   e   ������������������������       �                     @   E   ������������������������       �                      @f���  �       �                    �?�q�q�?             "@ v��  �       �                    �?�q�q�?             @    e   ������������������������       �                     �?*��  ������������������������       �                      @   e   �       �                 �UA@r�q��?             @       �       �                   @A@      �?             @    '   ������������������������       �                     �?    x   ������������������������       �                     @����  ������������������������       �                      @    "   �       �                 ���@�~�@
�?�            �x@    j   �       �                    7@�g�y��?             ?@    _   �       �                 03�@ףp=
�?             $@S��  ������������������������       �                     "@��  ������������������������       �                     �?    s   ������������������������       �                     5@��  �       
                ��Y7@�?��+�?�             w@   p   �       �                    /@����I�?�            �t@ ���  �       �                    $@      �?             8@   e   ������������������������       �        	             .@���  �       �                 �&�)@�q�q�?             "@    _   ������������������������       �                     @    e   �       �                    �?      �?             @ ���  ������������������������       �                      @   t   �       �                   �-@      �?              @    o   ������������������������       �                     �?�8��  ������������������������       �                     �?    m   �       �                    �?����Y��?�            s@    t   �       �                    �?���ȫ�?/            �T@    h   �       �                    �?�MI8d�?            �B@{��  �       �                    �?      �?             @@   o   ������������������������       �                     6@e   x   �       �                  S�-@z�G�z�?             $@    e   ������������������������       �                      @\и�  ������������������������       �                      @   t   �       �                 `�@1@z�G�z�?             @@��  ������������������������       �                     @        ������������������������       �                     �?`���  �       �                     @X�<ݚ�?            �F@׸�  �       �                  s@~�4_�g�?             F@    n   ������������������������       �                     @       �       �                   �3@      �?             D@ `��  ������������������������       �                     �?�и�  �       �                   �4@�99lMt�?            �C@ 3��  ������������������������       �                     @]   :   �       �                 ��/@b�2�tk�?             B@���  �       �                    �?�z�G��?             >@   m   �       �                   �5@�û��|�?             7@ ��  ������������������������       �                     �?    b   �       �                    �?���|���?             6@a��  �       �                   P&@�q�q�?             5@���  �       �                 �|�;@�z�G��?             4@       �       �                 pf�@�n_Y�K�?             *@ ���  ������������������������       �                      @�  �       �                 pf� @���!pc�?             &@b��  �       �                   �9@և���X�?             @:��  �       �                   �6@z�G�z�?             @    u   ������������������������       �                     �?"   "   ������������������������       �                     @MU��  ������������������������       �                      @�T��  ������������������������       �                     @       �       �                 ��� @؇���X�?             @   
   ������������������������       �                     @pY��  �       �                  SE"@      �?              @ Ը�  ������������������������       �                     �?����  ������������������������       �                     �?        ������������������������       �                     �?�t��  ������������������������       �                     �?f   r   ������������������������       �                     @�ĸ�  �       �                    �?r�q��?             @ |��  ������������������������       �                     �?�Ǹ�  ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?@�@+��?�            �k@    p   �       �                    �?�<ݚ�?             2@       �       �                   @@$�q-�?
             *@ o��  �       �                 �|�:@      �?             @ ��  ������������������������       �                      @�ո�  ������������������������       �      �?              @�o��  ������������������������       �                     "@        �       �                   �2@���Q��?             @ ���  ������������������������       �                      @8:��  ������������������������       �                     @bX��  �       �                    �?�M��?}            �i@ n��  �       �                    �?XB���?             =@��  ������������������������       �                     <@���  ������������������������       �                     �?    s   �       �                 �?�@h�V���?l             f@ i��  �       �                   �?@�k~X��?.             R@   -   ������������������������       �        %             L@<���  �       �                   @@@      �?	             0@    -   �       �                   �@      �?              @    -   ������������������������       �                     �?    -   ������������������������       �                     �?�ĸ�  ������������������������       �                     ,@i   c   �       �                   �1@�ջ����?>             Z@ j��  ������������������������       �                     (@-   -   �       	                   �?��H�?7             W@   -   �                          �?z�G�z�?2            @U@   -   �       �                 @3�@*�s���?1             U@ Ǹ�  �       �                   �?@      �?             ,@    m   �       �                   �9@�q�q�?             @       �       �                    �?      �?             @ ���  ������������������������       �                      @����  ������������������������       �                      @       ������������������������       �                      @   a   �       �                   �A@      �?              @ ��  ������������������������       ��q�q�?             @    l   ������������������������       ����Q��?             @        �       �                   �2@؇���X�?*            �Q@ ���  ������������������������       �                     @e   n   �       �                 ��) @pH����?)            �P@ ���  �       �                   �3@ 7���B�?             ;@ e��  ������������������������       �                     �?   _   ������������������������       �                     :@   g   �       �                   �9@R���Q�?             D@ ��  ������������������������       �                     1@   r   �                          (@��+7��?             7@R��  �                          ?@���Q��?             .@   r                          �|Y=@      �?              @    p   ������������������������       �                     @                              �̜!@���Q��?             @        ������������������������       �                     �?                              �|�=@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                              ��T?@��-�=��?            �C@       ������������������������       �                     9@                                 �?����X�?             ,@        ������������������������       �                     @                                 @���|���?             &@                                @���Q��?             $@                             ��p@@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �t�b�values�h*h-K ��h/��R�(KMKK��h]�BP        {@     Pq@     �`@      f@      ^@     �\@      2@      G@      1@      F@      *@      (@              @      *@      "@      @              $@      "@      @      @      @      @      �?               @      @              @       @              @      @              @      @              @       @      @                       @      @      @@              9@      @      @      �?      @      �?                      @      @      �?              �?      @              �?       @               @      �?             �Y@      Q@      1@      @              @      1@             @U@      P@     @T@     �D@      @@      ,@      ,@      (@              @      ,@      @              @      ,@      @      ,@      @      @               @      @      @      @              �?      @       @      @      �?      @      �?       @              �?      �?      �?                      �?       @                      �?      @                      �?      2@       @      (@              @       @              �?      @      �?      �?              @      �?              �?      @             �H@      ;@     �H@      6@      @      2@              "@      @      "@      @      @      �?      �?              �?      �?              @       @      @                       @       @      @       @       @               @       @                      @      E@      @     �A@      @      *@      @      *@       @      @              @       @      @              �?       @               @      �?                       @      6@              @                      @      @      7@      @      1@              @      @      (@      �?              @      (@              @      @      @       @              �?      @              @      �?      @              @      �?                      @      .@     �O@              1@      .@      G@      �?      >@      �?      @               @      �?      �?              �?      �?                      ;@      ,@      0@       @      *@       @      @      @      �?              �?      @              @      @              @      @                       @      @      @      �?       @      �?                       @      @      �?      @      �?              �?      @               @             �r@      Y@      >@      �?      "@      �?      "@                      �?      5@             �p@     �X@     @m@     �W@      @      5@              .@      @      @              @      @      �?       @              �?      �?      �?                      �?     �l@     �R@      ?@     �I@      @      ?@       @      >@              6@       @       @       @                       @      @      �?      @                      �?      9@      4@      9@      3@              @      9@      .@              �?      9@      ,@      @              6@      ,@      5@      "@      ,@      "@              �?      ,@       @      ,@      @      ,@      @       @      @               @       @      @      @      @      @      �?              �?      @                       @      @              @      �?      @              �?      �?              �?      �?                      �?              �?      @              �?      @      �?                      @              �?      i@      7@      ,@      @      (@      �?      @      �?       @              �?      �?      "@               @      @       @                      @     @g@      3@      <@      �?      <@                      �?     �c@      2@     �Q@      �?      L@              .@      �?      �?      �?              �?      �?              ,@             �U@      1@      (@             �R@      1@      Q@      1@     �P@      1@      @      @       @      @       @       @       @                       @               @      @      @       @      �?      @       @      N@      $@              @      N@      @      :@      �?              �?      :@              A@      @      1@              1@      @      "@      @       @      @              @       @      @              �?       @       @       @                       @      @               @              �?              @             �A@      @      9@              $@      @      @              @      @      @      @       @      @              @       @              @              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ/��hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtK�huh*h-K ��h/��R�(KK���h|�B�?                             @���*1�?�           8�@     �Y@                           @�7����?            �G@ o u r                             �?Pa�	�?            �@@ y��                             �?z�G�z�?             @    p y ������������������������       �                     �?       @������������������������       �                     @      9@������������������������       �                     <@      @       	                 ��T?@؇���X�?             ,@       @������������������������       �                      @0i�y�  
                           @�q�q�?             @i�y�  ������������������������       �                     @i�y�  ������������������������       �                      @0i�y�         z                     @��?a�?�           ��@ i�y�         !                    �?V$�݆��?�            �r@ i�y�                           0Cd=@Pns��ޭ?O            �`@ i�y�                            @E@$Q�q�?"            �O@i�y�                          ���*@p���?             I@                                `f�)@�IєX�?	             1@      ;@������������������������       �                     (@      "@                           :@z�G�z�?             @                                   5@      �?              @      @������������������������       �                     �?      @������������������������       �                     �?       @������������������������       �                     @       @������������������������       �                    �@@                                   �?�θ�?             *@     1@                        ���;@ףp=
�?             $@     (@������������������������       �                     "@      @������������������������       �                     �?                                   �?�q�q�?             @      G@������������������������       �                      @      �?������������������������       �                     �?      0@������������������������       �        -            �Q@      �?"       y                    �?4>���?t             e@       #       8                 `ff:@�{��?��?n            @d@        $       '                    5@ >�֕�?0            �Q@      �?%       &                   �2@      �?              @      �?������������������������       �                     �?        ������������������������       �                     �?      .@(       )                 �|Y=@ =[y��?.             Q@        ������������������������       �                     4@     �R@*       7                   �*@      �?#             H@     6@+       ,                 `f�)@ȵHPS!�?             :@     �?������������������������       �                     0@      3@-       .                 �|�=@�z�G��?             $@      ,@������������������������       �                     �?      "@/       4                   @D@�<ݚ�?             "@     @0       3                   �A@؇���X�?             @      @1       2                    @@�q�q�?             @       @������������������������       �                      @      �?������������������������       �                     �?      �?������������������������       �                     @      @5       6                   �G@      �?              @      �?������������������������       �                     �?        ������������������������       �                     �?      3@������������������������       �                     6@      2@9       V                    �?�)
;&��?>             W@      �?:       U                     �?�e����?            �C@     1@;       T                   �H@��J�fj�?            �B@     1@<       Q                   @C@�g�y��?             ?@       =       >                   �4@�û��|�?             7@      �?������������������������       �                     @      @?       P                 �̾w@�G�z��?             4@     @@       M                    �?ҳ�wY;�?             1@     @A       D                 �|�;@�q�q�?
             (@ ��  B       C                 Ȉ�P@�q�q�?             @     �?������������������������       �                      @      �?������������������������       �                     �?`���  E       L                   �A@�<ݚ�?             "@6��  F       K                 ��2>@�q�q�?             @        G       H                 `f&;@�q�q�?             @ ��  ������������������������       �                     �?       I       J                 ���<@      �?              @ ��  ������������������������       �                     �?�-��  ������������������������       �                     �?0��  ������������������������       �                     @�'��  ������������������������       �                     @        N       O                   �7@���Q��?             @ 4��  ������������������������       �                      @        ������������������������       �                     @���  ������������������������       �                     @p��  R       S                 ���X@      �?              @��  ������������������������       �                     @        ������������������������       �                     �?p��  ������������������������       �                     @����  ������������������������       �                      @p��  W       f                  i?@�c�����?"            �J@        X       e                   @>@p�ݯ��?             3@#��  Y       d                   �J@�t����?
             1@       Z       c                 `f�;@X�<ݚ�?             "@       [       ^                 �|�?@����X�?             @        \       ]                 �|�<@      �?              @  ��  ������������������������       �                     �?       ������������������������       �                     �?        _       `                   �C@z�G�z�?             @ ���  ������������������������       �                     @�*��  a       b                    H@      �?              @        ������������������������       �                     �?       ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @       ������������������������       �                      @pM��  g       x                     �?@�0�!��?             A@       h       i                   �A@�n`���?             ?@ ��  ������������������������       �                     "@�=��  j       w                    �?���!pc�?             6@���  k       v                    �?����X�?             5@���  l       m                   �B@�z�G��?             4@ ���  ������������������������       �                     @0��  n       u                 `f�K@@�0�!��?             1@       o       p                   �C@��S�ۿ?             .@��  ������������������������       �                     "@����  q       r                    �?r�q��?             @ @��  ������������������������       �                     @        s       t                  x#J@      �?              @        ������������������������       �                     �?       ������������������������       �                     �?���  ������������������������       �                      @        ������������������������       �                     �?p���  ������������������������       �                     �?0��  ������������������������       �                     @����  ������������������������       �                     @���  {       �                   �@@\�Yf�?�            �v@��  |       �                    �?�8a�ME�?�            �s@ ���  }       �                    �?@��Pl3�?<            @X@ ���  ~       �                    �?     ��?             @@F��         �                    �?�>4և��?             <@       �       �                    �?�IєX�?             1@ ��  ������������������������       �                      @       �       �                 �|�6@��S�ۿ?
             .@    p   ������������������������       �                     @    s   �       �                 ���@�8��8��?             (@    f   ������������������������       �                     �?        ������������������������       �                     &@       �       �                    �?���|���?             &@        �       �                   �,@z�G�z�?             @    n   ������������������������       �                     �?        ������������������������       �                     @    o   ������������������������       �                     @    t   ������������������������       �                     @        �       �                    �?&����?(            @P@       �       �                 03�-@>���Rp�?%             M@   s   �       �                    �?�LQ�1	�?             G@   S   �       �                    �?8�Z$���?             :@       �       �                 ���@r�q��?             8@    T   ������������������������       �                     "@   t   �       �                   @@������?             .@   y   �       �                   �5@�q�q�?             "@    t   ������������������������       �                     �?        �       �                 �|=@      �?              @    ,   ������������������������       �                      @    y   �       �                 �|�=@�q�q�?             @       ������������������������       �      �?             @    o   ������������������������       �                      @       �       �                 �|Y=@r�q��?             @    n   ������������������������       �                     �?   m   ������������������������       �                     @    i   ������������������������       �                      @        �       �                 �|Y;@ףp=
�?             4@    e   ������������������������       �                     �?    
   �       �                  s�@�KM�]�?             3@        ������������������������       �                     @   _   �       �                    �?؇���X�?
             ,@       ������������������������       �8�Z$���?	             *@       ������������������������       �                     �?   i   �       �                 ��.@�q�q�?             (@    y   ������������������������       �                     @       �       �                 ��$1@և���X�?             @    n   ������������������������       �                     @    o   �       �                   �2@      �?             @    b   ������������������������       �                     �?       ������������������������       �                     @       ������������������������       �                     @   t   �       �                    �?�nYU}�?�             k@       �       �                    @�C�F��?o            �e@       �       �                 �|�=@�R����?n            �e@   l   �       �                    �?*~k���?b            �b@    .   �       �                  s@�eP*L��?             6@    n   ������������������������       �                     @       �       �                    4@�q�q�?             2@        �       �                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?    v   �       �                 �|�;@d}h���?
             ,@       �       �                 pff@ףp=
�?             $@        �       �                   �7@      �?              @        ������������������������       �                     �?    e   ������������������������       �                     �?    a   ������������������������       �                      @        �       �                    �?      �?             @   v   ������������������������       �                      @       ������������������������       �                      @       �       �                    �?x�]AgȽ?T             `@   F   �       �                    �?`Jj��?R             _@       �       �                 ���@�IєX�?N            �]@ K@lt ��       �                   �5@����X�?             @    
   ������������������������       �                     @        �       �                 �&b@      �?             @   ,   ������������������������       �                      @G   r   ������������������������       �                      @        �       �                   �0@���>4ֵ?I             \@    r   �       �                 pFD!@      �?             @    t   ������������������������       �      �?              @   c   ������������������������       �                      @        �       �                 @3�!@ 7���B�?E             [@   i   �       �                 @3�@������?6            �T@   p   �       �                 �?$@���J��?!            �I@    )   �       �                 ��@���N8�?             5@       ������������������������       �        	             1@    l   �       �                 �|Y8@      �?             @        ������������������������       �                     �?   t   ������������������������       ��q�q�?             @   a   ������������������������       �                     >@        �       �                 pf� @��a�n`�?             ?@   p   �       �                   �4@�8��8��?             8@        �       �                   �2@����X�?             @        ������������������������       �                      @   t   �       �                 0S5 @���Q��?             @   e   ������������������������       ��q�q�?             @       ������������������������       �                      @       ������������������������       �                     1@       �       �                    8@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?    t   ������������������������       �                     :@       �       �                 �Y�@z�G�z�?             @        ������������������������       �                      @       �       �                 pF�+@�q�q�?             @        ������������������������       �                     �?    e   ������������������������       �                      @   n   ������������������������       �                     @    x   �       �                   @@@8�A�0��?             6@   i   �       �                    �?      �?
             2@       �       �                    �?     ��?	             0@    #   ������������������������       �                     @   .   �       �                   �?@��
ц��?             *@    t   ������������������������       �                     @    t   �       �                 d�6@@���Q��?             $@       �       �                 ��I @և���X�?             @       �       �                 P�@      �?             @    a   ������������������������       �                      @    r   ������������������������       �      �?              @       ������������������������       �                     @       ������������������������       �                     @       ������������������������       �                      @    _   ������������������������       �                     @       ������������������������       �                      @        �       �                 �̜2@d}h���?             E@        �       �                    <@�	j*D�?             *@       �       �                 P�@"pc�
�?             &@    s   ������������������������       �                      @    a   ������������������������       �                     "@   r   ������������������������       �                      @        ������������������������       �                     =@        ������������������������       �                     H@        �t�bh�h*h-K ��h/��R�(KK�KK��h]�B�       �{@     �p@      *@      A@      �?      @@      �?      @      �?                      @              <@      (@       @       @              @       @      @                       @     �z@     �m@     �a@     @d@      @      `@      @     �M@      �?     �H@      �?      0@              (@      �?      @      �?      �?              �?      �?                      @             �@@      @      $@      �?      "@              "@      �?               @      �?       @                      �?             �Q@      a@     �@@      `@     �@@     �P@      @      �?      �?      �?                      �?     @P@      @      4@             �F@      @      7@      @      0@              @      @              �?      @       @      @      �?       @      �?       @                      �?      @              �?      �?              �?      �?              6@             �O@      =@      7@      0@      5@      0@      .@      0@      ,@      "@      @              &@      "@      &@      @       @      @      �?       @               @      �?              @       @      @       @      �?       @              �?      �?      �?      �?                      �?      @              @              @       @               @      @                      @      �?      @              @      �?              @               @              D@      *@      (@      @      (@      @      @      @       @      @      �?      �?              �?      �?              �?      @              @      �?      �?      �?                      �?       @               @                       @      <@      @      9@      @      "@              0@      @      .@      @      ,@      @              @      ,@      @      ,@      �?      "@              @      �?      @              �?      �?      �?                      �?               @      �?              �?              @              @             �q@     �R@     �m@     �R@      N@     �B@      "@      7@      @      7@      �?      0@               @      �?      ,@              @      �?      &@      �?                      &@      @      @      @      �?              �?      @                      @      @             �I@      ,@      F@      ,@      D@      @      6@      @      4@      @      "@              &@      @      @      @              �?      @       @       @              @       @       @       @       @              @      �?              �?      @               @              2@       @      �?              1@       @      @              (@       @      &@       @      �?              @       @              @      @      @      @              �?      @      �?                      @      @             `f@      C@     @b@      =@     @b@      ;@     �`@      2@      (@      $@              @      (@      @      �?      @              @      �?              &@      @      "@      �?      �?      �?              �?      �?               @               @       @       @                       @     @^@       @      ]@       @      \@      @      @       @      @               @       @       @                       @     �Z@      @      @      �?      �?      �?       @              Z@      @     �S@      @      I@      �?      4@      �?      1@              @      �?      �?               @      �?      >@              <@      @      6@       @      @       @       @              @       @      �?       @       @              1@              @      �?      @                      �?      :@              @      �?       @               @      �?              �?       @              @              *@      "@      "@      "@      @      "@              @      @      @      @              @      @      @      @      �?      @               @      �?      �?      @                      @       @              @                       @     �@@      "@      @      "@       @      "@       @                      "@       @              =@              H@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJu�7hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B�F         D                    �?���Yb�?�           8�@     �Y@       )                    �?&ջ�{��?]            @b@���                             �?JJ����?;            �W@ 6��                             �?��hJ,�?             A@3��  ������������������������       �                     ;@      @                        �ܙH@����X�?             @     @������������������������       �                     @      "@������������������������       �                      @      �?	       
                   �2@      �?'             N@      @������������������������       �                     @     �D@                             @����>4�?$             L@      @                          @B@�ՙ/�?             5@                               ���<@      �?             0@       @������������������������       �                     @      �?                           �?�n_Y�K�?	             *@     �?                        03SA@���Q��?             $@        ������������������������       �                     @                                @�6M@և���X�?             @      �?������������������������       �                     @                                X�,@@      �?             @                               �|Y<@      �?              @        ������������������������       �                     �?      @������������������������       �                     �?      �?������������������������       �                      @      @                        �nc@�q�q�?             @        ������������������������       �                     �?      @                        �̾w@      �?              @      @������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @               "                 �|Y=@�#-���?            �A@     �R@        !                   @@z�G�z�?             $@     0@������������������������       �                      @Ɂ��  ������������������������       �                      @�8��  #       $                 ���@`2U0*��?             9@ ���  ������������������������       �                     &@0���  %       (                 �|�=@@4և���?
             ,@���  &       '                   @@      �?              @>��  ������������������������       �r�q��?             @0��  ������������������������       �                      @p��  ������������������������       �                     @0��  *       3                     @R�}e�.�?"             J@��  +       ,                    �?z�G�z�?             >@��  ������������������������       �                     4@0���  -       2                    �?���Q��?             $@     �?.       1                     �?�q�q�?             @���  /       0                 �U�X@z�G�z�?             @��  ������������������������       �                     @0���  ������������������������       �                     �?(N��  ������������������������       �                     �?0���  ������������������������       �                     @      @4       =                    �?���|���?
             6@ ���  5       <                    �?և���X�?             ,@���  6       9                    �?�eP*L��?             &@ ���  7       8                   �-@և���X�?             @ ���  ������������������������       �                     @���  ������������������������       �                     @p���  :       ;                 �|Y3@      �?             @ ���  ������������������������       �                     @0��  ������������������������       �                     �?0<��  ������������������������       �                     @����  >       C                 03�-@      �?              @���  ?       B                    �?�q�q�?             @b��  @       A                 �&�)@      �?              @ ��  ������������������������       �                     �? ��  ������������������������       �                     �?     �?������������������������       �                     �?      �?������������������������       �                     @`���  E                       `f�S@��f
a�?r           ��@6��  F       �                 `f�$@�K�7���?]           Ȁ@        G       \                    �?��1��?�            �n@ ��  H       S                   �6@�g�y��?             ?@        I       R                    �?r�q��?
             (@��  J       O                    �?�<ݚ�?             "@-��  K       L                    �?؇���X�?             @ ��  ������������������������       �                      @�'��  M       N                   �3@z�G�z�?             @        ������������������������       �                     �? 4��  ������������������������       �                     @        P       Q                    4@      �?              @ ��  ������������������������       �                     �?p��  ������������������������       �                     �?��  ������������������������       �                     @        T       Y                 ��@�d�����?             3@ ��  U       V                 ���@�q�q�?             @ ���  ������������������������       �                     �?p��  W       X                    �?z�G�z�?             @       ������������������������       �                     @#��  ������������������������       �                     �?       Z       [                    �?$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@  ��  ]       b                   �0@d��]a��?�            �j@        ^       _                 pf�@���!pc�?             &@        ������������������������       �                     @ ���  `       a                 pFD!@և���X�?             @ *��  ������������������������       �                     @        ������������������������       �                     @       c       l                    �?����p�?�            �i@        d       e                 ���@�>4և��?             <@        ������������������������       �                      @       f       g                 �|Y=@      �?
             4@ M��  ������������������������       �                     @       h       k                 X��A@�t����?	             1@��  i       j                    �?؇���X�?             ,@=��  ������������������������       �8�Z$���?             *@���  ������������������������       �                     �?���  ������������������������       �                     @ ���  m       �                 �|�=@����!p�?u             f@��  n       {                 �?$@ ,V�ނ�?V            �_@        o       x                 ���@�L���?            �B@��  p       q                     @�g�y��?             ?@ ���  ������������������������       �                     "@ @��  r       s                  Md@���7�?             6@        ������������������������       �                     &@        t       u                    7@�C��2(�?             &@        ������������������������       �                     @���  v       w                   �8@r�q��?             @        ������������������������       �                     �?p���  ������������������������       �                     @0��  y       z                 �|�;@�q�q�?             @ ���  ������������������������       �                     @���  ������������������������       ��q�q�?             @��  |       �                    �?�x�E~�?;            @V@���  }       �                    �?`���i��?:             V@���  ~                        @3�@�D�e���?8            @U@ F��  ������������������������       �                    �C@       �       �                   �;@�nkK�?             G@��  �       �                   �9@�>����?             ;@��z�  �       �                   �3@ ��WV�?             :@ Wz�  �       �                   �2@�C��2(�?             &@ ��z�  ������������������������       �                     @ Xz�  �       �                 0S5 @؇���X�?             @ TMy� �������������������������       �      �?              @ �z�  ������������������������       �                     @��z�  ������������������������       �        	             .@Sz�  ������������������������       �                     �? Uz�  ������������������������       �                     3@Qz�  ������������������������       �                     @ Uz�  ������������������������       �                     �?pVz�  �       �                   @@@ףp=
�?             I@ Uz�  �       �                 �?�@�	j*D�?             *@ Wz�  ������������������������       �                     @�z�  �       �                    ?@X�<ݚ�?             "@ �z�  �       �                 �̌!@      �?              @ �z�  ������������������������       �                     �? ��z�  ������������������������       �                     �? �z�  �       �                 ��I @և���X�?             @�z�  ������������������������       ����Q��?             @�z�  ������������������������       �                      @ �z�  �       �                      @�?�|�?            �B@ ��z�  ������������������������       �                     @ ��z�  �       �                   �C@г�wY;�?             A@�z�  �       �                   @C@�IєX�?             1@�z�  ������������������������       �        
             .@�z�  ������������������������       �      �?              @l�y�  ������������������������       �        	             1@Uz�  �       �                    �?��c���?�            0r@ Qz�  �       �                    �?ڷv���?I            �\@ Wz�  �       �                    �?Hm_!'1�?            �H@ �z�  ������������������������       �                     �? �z�  �       �                    �?      �?             H@�z�  �       �                     @ �Cc}�?             <@��z�  �       �                     �?$�q-�?             :@ �z�  ������������������������       �                     @��z�  �       �                   �A@�C��2(�?             6@�z�  �       �                   �9@�IєX�?
             1@ Tz�  �       �                   �'@؇���X�?             @ Vz�  ������������������������       �                     @���z�  �       �                   �3@      �?              @ ��z�  ������������������������       �                     �?�z�  ������������������������       �                     �? �z�  ������������������������       �                     $@ Rz�  �       �                   �D@z�G�z�?             @ Uz�  ������������������������       �                     �? Wz�  ������������������������       �                     @ �z�  �       �                 ��&@      �?              @ ��z�  ������������������������       �                     �?�z�  ������������������������       �                     �? Tz�  ������������������������       �                     4@ Vz�  �       �                     @8�A�0��?*            �P@ ��z�  �       �                     �?�}�+r��?             3@ Uz�  ������������������������       �                     @Wz�  �       �                    �?��S�ۿ?             .@ j�y�  �       �                    B@      �?             @��z�  ������������������������       �                     @��z�  ������������������������       �                     �?�z�  ������������������������       �        	             &@Vz�  �       �                    �?��k=.��?            �G@ Wz�  ������������������������       �                      @ �z�  �       �                   @1@���V��?            �F@ Qz�  �       �                    �?���|���?             &@Wz�  �       �                    D@����X�?             @�z�  �       �                 �|�;@      �?             @ �z�  ������������������������       �                      @�z�  ������������������������       �                      @ �z�  ������������������������       �                     @ �z�  �       �                    0@      �?             @ Uz�  ������������������������       �                      @ l�y�  ������������������������       �                      @Wz�  �       �                    @l��\��?             A@ Wz�  �       �                    @����X�?             @Sz�  ������������������������       �                     @ �z�  ������������������������       �                      @ �z�  �       �                    @ 7���B�?             ;@Wz�  ������������������������       �                     7@��z�  �       �                   @D@      �?             @ �z�  ������������������������       �                     �?�z�  ������������������������       �                     @ �z�  �                          �?��|���?t             f@Tz�  �       �                    �?H%u��?T            @_@ Vz�  �       �                    �?      �?              @��z�  ������������������������       �                     @�z�  ������������������������       �                     �?��z�  �       �                 `fF:@�S#א��?N            @]@�z�  �       �                    4@����p�?+             Q@ �z�  �       �                    &@�<ݚ�?             "@ ��z�  ������������������������       �                      @Wz�  ������������������������       �                     @�z�  �       �                     @����˵�?$            �M@��z�  �       �                   �*@���.�6�?             G@Uz�  �       �                 `f�)@ܷ��?��?             =@ Wz�  ������������������������       �                     @ �z�  �       �                   �A@�LQ�1	�?             7@�z�  �       �                    @@d}h���?             ,@�z�  ������������������������       �                      @ m�y�  ������������������������       �      �?             @ �z�  ������������������������       �                     "@�z�  ������������������������       �                     1@ �z�  ������������������������       �                     *@�z�  �                         �Q@Jm_!'1�?#            �H@i�y�  �                          �?r�q��?"             H@   s   �                             @t/*�?!            �G@   #   �       �                   �;@"pc�
�?             F@    k   �       �                    �?�q�q�?             @    g   ������������������������       �                     �?   i   �       �                    7@      �?              @    b   ������������������������       �                     �?        ������������������������       �                     �?   p   �       �                   �>@�p ��?            �D@    t   �       �                    K@     ��?             0@   f   �       �                   `G@�eP*L��?             &@   g   �       �                   @>@      �?              @   _   �       �                 `f�;@؇���X�?             @   l   �       �                 �|�<@      �?             @        ������������������������       �                     �?    s   ������������������������       �                     @    a   ������������������������       �                     @        ������������������������       �                     �?   a   ������������������������       �                     @       ������������������������       �                     @       �       �                  x#J@`2U0*��?             9@   a   ������������������������       �                     1@   f   �       �                 `�iJ@      �?              @    e   ������������������������       �                     �?       ������������������������       �                     @    t   ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?                                 �?��[�8��?             �I@                                +@J�8���?             =@        ������������������������       �                     $@        ������������������������       �                     3@                                 @���7�?             6@       	      
                   �?      �?
             0@       ������������������������       �                     *@                                 @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                 �?�>4և��?             <@                                M@H%u��?             9@                              �k@�8��8��?             8@                               @E@�nkK�?             7@       ������������������������       �                     3@                                 �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?                                 @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �t�bh�h*h-K ��h/��R�(KMKK��h]�B�       �}@     �m@      P@     �T@      I@      F@      @      =@              ;@      @       @      @                       @     �F@      .@              @     �F@      &@      *@       @       @       @      @              @       @      @      @              @      @      @      @              �?      @      �?      �?              �?      �?                       @      �?       @              �?      �?      �?      �?                      �?      @              @@      @       @       @       @                       @      8@      �?      &@              *@      �?      @      �?      @      �?       @              @              ,@      C@      @      8@              4@      @      @       @      @      �?      @              @      �?              �?              @               @      ,@      @       @      @      @      @      @      @                      @      @      �?      @                      �?              @       @      @       @      �?      �?      �?              �?      �?              �?                      @     �y@     @c@     `y@     ``@     �j@     �@@      0@      .@       @      $@       @      @      �?      @               @      �?      @      �?                      @      �?      �?              �?      �?                      @      ,@      @       @      @      �?              �?      @              @      �?              (@      �?              �?      (@             �h@      2@       @      @      @              @      @              @      @             �g@      .@      7@      @       @              .@      @              @      .@       @      (@       @      &@       @      �?              @             �d@      $@     @^@      @      A@      @      >@      �?      "@              5@      �?      &@              $@      �?      @              @      �?              �?      @              @       @      @              �?       @     �U@       @     �U@       @     �T@       @     �C@              F@       @      9@       @      9@      �?      $@      �?      @              @      �?      �?      �?      @              .@                      �?      3@              @              �?             �F@      @      "@      @      @              @      @      �?      �?      �?                      �?      @      @       @      @       @              B@      �?      @             �@@      �?      0@      �?      .@              �?      �?      1@              h@     �X@     �E@      R@      @     �F@      �?              @     �F@      @      9@       @      8@              @       @      4@      �?      0@      �?      @              @      �?      �?      �?                      �?              $@      �?      @      �?                      @      �?      �?      �?                      �?              4@     �C@      ;@      �?      2@              @      �?      ,@      �?      @              @      �?                      &@      C@      "@               @      C@      @      @      @      @       @       @       @       @                       @      @               @       @               @       @              ?@      @      @       @      @                       @      :@      �?      7@              @      �?              �?      @             �b@      :@     �[@      .@      @      �?      @                      �?     �Y@      ,@     �O@      @      @       @               @      @              L@      @     �E@      @      :@      @      @              4@      @      &@      @       @              @      @      "@              1@              *@              D@      "@      D@       @     �C@       @      B@       @      �?       @              �?      �?      �?      �?                      �?     �A@      @      &@      @      @      @      @       @      @      �?      @      �?              �?      @              @                      �?              @      @              8@      �?      1@              @      �?              �?      @              @              �?                      �?      D@      &@      3@      $@              $@      3@              5@      �?      .@      �?      *@               @      �?       @                      �?      @              @      7@      @      6@       @      6@      �?      6@              3@      �?      @              @      �?              �?              �?               @      �?       @                      �?�t�bub�$>     hhubh)��}�(hhhhhNhKhKhG        hh&hNhJ��!XhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM	huh*h-K ��h/��R�(KM	��h|�B@B         l                 ��%@�*���?�           8�@      @                           /@,PY��?�             v@ ���  ������������������������       �                     @      =@                        ���@j�q����?�            �u@      *@������������������������       �                    �E@      @       3                 P�*@�A��t��?�            0s@       @       2                 �|Y>@J��D��?A             [@              1                    �?���Q �?8            �X@      @	       
                 ��@r�qG�?7             X@        ������������������������       �                     �?                                   �?�|R���?6            �W@                                  �3@���B���?             :@                                �?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �?�LQ�1	�?             7@                                  8@�C��2(�?             6@        ������������������������       �                     "@      ;@                        ��@8�Z$���?	             *@     "@                        ���@�C��2(�?             &@                                   �?�q�q�?             @      @������������������������       �                      @      @������������������������       �                     �?       @������������������������       �                      @       @                           @      �?              @        ������������������������       �                     �?     1@������������������������       �                     �?     (@������������������������       �                     �?      @       $                   �<@�㙢�c�?&            @Q@               #                   �6@�C��2(�?            �@@     G@                           �3@�S����?
             3@      �?������������������������       �                      @      0@!       "                    �?���!pc�?             &@      @������������������������       �                     @      @������������������������       �                      @        ������������������������       �                     ,@      @%       .                    �?      �?             B@       &       '                 ���@z�G�z�?             9@        ������������������������       �                      @     @(       )                 �|Y=@�t����?             1@        ������������������������       �                     �?     @*       +                 ���@      �?
             0@       @������������������������       ����Q��?             @        ,       -                 �Y�@�C��2(�?             &@       @������������������������       �                     @       @������������������������       �      �?              @    �A@/       0                 ��,@���|���?             &@     :@������������������������       �                     @       @������������������������       ��q�q�?             @       ������������������������       �                      @      "@������������������������       �        	             $@       @4       i                    �?ȭ^���?x            �h@       5       <                 �?�@��ɉ�?v            `h@      @6       ;                 �̌@�L#���?)            �P@      &@7       8                 �|Y=@���y4F�?             3@      @������������������������       �        
             *@        9       :                 ��]@�q�q�?             @       @������������������������       �                      @        ������������������������       �                     @      @������������������������       �                     H@      @=       B                     @     ��?M             `@      �?>       A                   �J@�+e�X�?             9@       ?       @                    �?�����?             3@      @������������������������       �                     @      @������������������������       �                     *@       @������������������������       �                     @        C       N                 @3�@�v�G���??            �Y@        D       G                    �?      �?             0@      @E       F                   �9@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        H       I                    :@���|���?             &@        ������������������������       �                     @        J       K                   �?@և���X�?             @        ������������������������       �                     �?        L       M                   �A@      �?             @        ������������������������       �      �?              @        ������������������������       �      �?             @        O       V                   �:@�=C|F�?4            �U@        P       U                   �3@`Ӹ����?            �F@        Q       T                 0S5 @�����?
             5@        R       S                   �1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     2@        ������������������������       �                     8@        W       X                   �;@d}h���?             E@        ������������������������       �                     @        Y       h                   �?@8�Z$���?            �C@       Z       [                 ��) @      �?             8@       ������������������������       �        	             &@        \       ]                   �<@��
ц��?             *@        ������������������������       �                     @        ^       c                 P�*"@���Q��?             $@        _       `                 pf� @z�G�z�?             @        ������������������������       �                      @        a       b                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        d       e                 ���"@���Q��?             @        ������������������������       �                      @        f       g                 �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             .@        j       k                   �#@      �?             @        ������������������������       �                      @        ������������������������       �                      @        m       �                  x#J@��d���?�            Pv@       n       �                    �?~���n��?�            Pp@        o       �                    @t�I��n�?R            @]@       p       u                    @f�����?N            �[@        q       r                    @�}�+r��?             3@       ������������������������       �        
             0@        s       t                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        v       �                     @ �&�T�?B             W@       w       �                   �H@�j��b�?(            �M@       x       �                    �?,�+�C�?%            �K@       y       z                     �?<���D�?            �@@        ������������������������       �                     @        {       �                   �7@8�Z$���?             :@       |       �                    �?������?             .@       }       �                    :@d}h���?             ,@        ~                           �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?ףp=
�?	             $@ ��z�  ������������������������       �                     �? Wz�  �       �                   �*@�����H�?             "@��z�  �       �                 `f�)@؇���X�?             @ Xz�  ������������������������       �                     �? TMy� ��       �                   �B@r�q��?             @�z�  ������������������������       �                     @��z�  ������������������������       �                     �?Sz�  ������������������������       �                      @ Uz�  ������������������������       �                     �?Qz�  ������������������������       �                     &@ Uz�  ������������������������       �                     6@pVz�  �       �                 03�9@      �?             @Uz�  ������������������������       �                      @ Wz�  ������������������������       �                      @�z�  �       �                    �?4���C�?            �@@�z�  �       �                 ��.@\X��t�?             7@�z�  �       �                    �?�	j*D�?
             *@ ��z�  �       �                 �|Y6@և���X�?             @�z�  �       �                   �,@      �?             @ �z�  ������������������������       �                      @�z�  �       �                   �-@      �?              @ �z�  ������������������������       �                     �? ��z�  ������������������������       �                     �? ��z�  ������������������������       �                     @�z�  �       �                   �*@r�q��?             @ �z�  ������������������������       �                     �?�z�  ������������������������       �                     @l�y�  �       �                    �?ףp=
�?             $@ Uz�  ������������������������       �                     @ Qz�  �       �                 �|Y>@r�q��?             @ Wz�  ������������������������       �                     @ �z�  �       �                 03C3@      �?              @ �z�  ������������������������       �                     �?�z�  ������������������������       �                     �?��z�  �       �                 ���0@ףp=
�?             $@ �z�  ������������������������       �                     �?��z�  ������������������������       �                     "@�z�  ������������������������       �                     @ Tz�  �       �                    @�q�q�?g             b@Vz�  �       �                    !@�θ�?^            @`@ ��z�  ������������������������       �                     $@ ��z�  �       �                 �&@r�q��?W             ^@ �z�  ������������������������       �                     �? �z�  �       �                     �?�?��,�?V            �]@ Rz�  �       �                 ��";@���j��?             G@ Uz�  �       �                 ��$:@և���X�?
             ,@ Wz�  ������������������������       �                     @ �z�  �       �                   �J@���!pc�?             &@��z�  �       �                   @G@�����H�?             "@�z�  �       �                    D@z�G�z�?             @ Tz�  ������������������������       �                      @ Vz�  ������������������������       ��q�q�?             @ ��z�  ������������������������       �                     @ Uz�  ������������������������       �                      @Wz�  �       �                    �?     ��?             @@j�y�  �       �                 ���=@�����?             5@ ��z�  ������������������������       �                     $@��z�  �       �                 p�i@@"pc�
�?             &@ �z�  �       �                 �|�;@�q�q�?             @ Vz�  ������������������������       �                     �? Wz�  �       �                  �>@      �?              @ �z�  ������������������������       �                     �? Qz�  ������������������������       �                     �?Wz�  ������������������������       �                      @�z�  �       �                   �<@���!pc�?	             &@ �z�  ������������������������       �                      @�z�  �       �                 �|Y>@�����H�?             "@ �z�  �       �                 �|Y=@      �?             @ �z�  ������������������������       �                     �? Uz�  �       �                   �>@�q�q�?             @ l�y�  ������������������������       �                     �?Wz�  ������������������������       �                      @ Wz�  ������������������������       �                     @Sz�  �       �                   �*@�F��O�?8            @R@ �z�  �       �                   �@@�㙢�c�?             7@�z�  ������������������������       �        
             (@Wz�  �       �                   �)@���|���?	             &@ �z�  ������������������������       �                      @ �z�  �       �                   �A@X�<ݚ�?             "@ �z�  ������������������������       �      �?             @ �z�  �       �                   @D@z�G�z�?             @ Tz�  ������������������������       �                      @ Vz�  �       �                    G@�q�q�?             @ ��z�  ������������������������       �                     �?�z�  ������������������������       �                      @��z�  �       �                    �?`2U0*��?%             I@�z�  �       �                 ��.@`Ql�R�?"            �G@ �z�  �       �                     @$�q-�?
             *@ ��z�  ������������������������       �                     @Wz�  �       �                    �?r�q��?             @�z�  ������������������������       �                     @��z�  �       �                    �?      �?              @ Uz�  ������������������������       �                     �? Wz�  ������������������������       �                     �? �z�  ������������������������       �                     A@�z�  �       �                    �?�q�q�?             @ �z�  ������������������������       �                     �? m�y�  ������������������������       �                      @ �z�  ������������������������       �        	             ,@�z�  �                          @     ��?B             X@�z�  �       �                    �?�n`���??            @W@�z�  �       �                   �5@f>�cQ�?-            �N@ i�y�  �       �                    �?X�<ݚ�?             "@    s   ������������������������       �                     @   #   ������������������������       �                     @    k   �       �                    �?$�q-�?'             J@   g   �       �                      @�IєX�?&            �I@   i   �       �                   �B@ �q�q�?#             H@   b   �       �                    �?�IєX�?             A@       ������������������������       �                     <@   p   �       �                    �?�q�q�?             @   t   �       �                 X�,@@      �?             @   f   �       �                 p"�b@      �?              @    g   ������������������������       �                     �?   _   ������������������������       �                     �?   l   ������������������������       �                      @        �       �                    �?      �?              @    s   ������������������������       �                     �?    a   ������������������������       �                     �?        ������������������������       �        
             ,@   a   �       �                 �|�;@�q�q�?             @        ������������������������       �                     �?       �       �                 �|�>@      �?              @    a   ������������������������       �                     �?   f   ������������������������       �                     �?    e   ������������������������       �                     �?                                �7@     ��?             @@    t                            �?�C��2(�?             &@                                �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                 �?�ՙ/�?             5@       ������������������������       �                     *@        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h*h-K ��h/��R�(KM	KK��h]�B�       `|@     p@     �q@     �P@              @     �q@     �O@     �E@             �n@     �O@     �R@      A@      P@      A@      O@      A@              �?      O@     �@@      @      5@       @      �?              �?       @              @      4@       @      4@              "@       @      &@      �?      $@      �?       @               @      �?                       @      �?      �?      �?                      �?      �?             �L@      (@      >@      @      0@      @       @               @      @              @       @              ,@              ;@      "@      4@      @       @              (@      @              �?      (@      @       @      @      $@      �?      @              @      �?      @      @      @               @      @       @              $@             @e@      =@      e@      ;@     �O@      @      .@      @      *@               @      @       @                      @      H@             @Z@      7@      3@      @      *@      @              @      *@              @             �U@      1@      $@      @      @       @      @                       @      @      @      @              @      @              �?      @      @      �?      �?       @       @      S@      &@     �E@       @      3@       @      �?       @      �?                       @      2@              8@             �@@      "@              @     �@@      @      2@      @      &@              @      @      @              @      @      �?      @               @      �?       @               @      �?              @       @       @              �?       @               @      �?              .@               @       @               @       @             �d@     �g@     @b@     �\@      @@     @U@      :@     @U@      �?      2@              0@      �?       @      �?                       @      9@     �P@      @     �J@      @     �I@      @      =@              @      @      6@      @      &@      @      &@       @       @               @       @              �?      "@              �?      �?       @      �?      @              �?      �?      @              @      �?                       @      �?                      &@              6@       @       @               @       @              3@      ,@      $@      *@      "@      @      @      @      �?      @               @      �?      �?      �?                      �?      @              @      �?              �?      @              �?      "@              @      �?      @              @      �?      �?      �?                      �?      "@      �?              �?      "@              @             �\@      >@      Y@      >@              $@      Y@      4@              �?      Y@      3@     �@@      *@      @       @      @              @       @      �?       @      �?      @               @      �?       @              @       @              ;@      @      3@       @      $@              "@       @      �?       @              �?      �?      �?      �?                      �?       @               @      @               @       @      �?      @      �?      �?               @      �?              �?       @              @             �P@      @      3@      @      (@              @      @       @              @      @      �?      @      @      �?       @               @      �?              �?       @              H@       @      G@      �?      (@      �?      @              @      �?      @              �?      �?      �?                      �?      A@               @      �?              �?       @              ,@              5@     �R@      2@     �R@      "@      J@      @      @              @      @              @      H@      @      H@       @      G@       @      @@              <@       @      @      �?      @      �?      �?              �?      �?                       @      �?      �?              �?      �?                      ,@      �?       @              �?      �?      �?      �?                      �?      �?              "@      7@      �?      $@      �?      @      �?                      @              @       @      *@              *@       @              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJC�NhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM	huh*h-K ��h/��R�(KM	��h|�B@B         p                     @���%&�?�           8�@      @       '                 �|Y=@N�ec�?�            ps@ paramet       
                 ��*@"��$�?G            �[@      @       	                    �?      �?             8@       @                           �?"pc�
�?             &@     $@                        `f�)@�<ݚ�?             "@      @������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        
             *@               "                 `fmj@�N��D�?6            �U@                                  �?���(\��?2             T@                                  6@�C��2(�?)            �P@                                   9@���|���?             &@       ������������������������       �                     @                                   �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @      ;@                           �?h㱪��?#            �K@     "@������������������������       �                    �B@                                    �?�����H�?
             2@     @                           5@��S�ۿ?             .@      @������������������������       �                     �?       @������������������������       �                     ,@       @                           �?�q�q�?             @        ������������������������       �                     �?     1@������������������������       �                      @     (@                           �?d}h���?	             ,@     @                            �?�����H�?             "@        ������������������������       �                     �?     G@������������������������       �                      @      �?        !                    �?���Q��?             @     0@������������������������       �                     @      @������������������������       �                      @      @#       &                 0U�o@և���X�?             @       $       %                    5@z�G�z�?             @      @������������������������       �                     �?       ������������������������       �                     @        ������������������������       �                      @     @(       9                    �?4��@���?�             i@        )       ,                    �?�nkK�?1            @Q@      @*       +                 03�=@`2U0*��?             9@       @������������������������       �                     �?        ������������������������       �                     8@       @-       6                    L@���7�?             F@      @.       /                   �B@��Y��]�?            �D@    �A@������������������������       �                     8@     :@0       5                    -@�IєX�?             1@       @1       2                   �'@�q�q�?             @        ������������������������       �                     �?      "@3       4                    D@      �?              @       @������������������������       �                     �?       ������������������������       �                     �?      @������������������������       �        	             ,@      &@7       8                   �L@�q�q�?             @       @������������������������       �                     �?        ������������������������       �                      @       @:       o                   �J@��ׂ�?Z            ``@       ;       n                 p�w@������?F            @Z@     @<       a                   �G@��z6��?D             Y@     @=       >                   �)@� ���?6            @S@      �?������������������������       �        	             ,@       ?       `                   �F@��s����?-            �O@     @@       [                    �?�T`�[k�?(            �J@     @A       L                    �?��Q���?             D@      &@B       K                    �?     ��?
             0@     �?C       J                    C@�q�q�?	             .@       D       I                 ��2>@����X�?             ,@      6@E       H                 ���<@      �?              @     @F       G                 ��";@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        M       Z                    �?      �?             8@       N       W                   @D@���!pc�?             6@       O       V                 `f�<@@�0�!��?             1@       P       U                 `fF:@���!pc�?             &@       Q       T                 `fv3@z�G�z�?             $@       R       S                 �|�=@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        X       Y                     �?���Q��?             @        ������������������������       �      �?              @        ������������������������       ��q�q�?             @        ������������������������       �                      @        \       ]                   �B@$�q-�?             *@        ������������������������       �                     @        ^       _                 03�U@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        b       c                 `f4@
;&����?             7@        ������������������������       �                     @        d       i                    �?     ��?	             0@        e       f                    �?�q�q�?             @        ������������������������       �                      @        g       h                 ���X@      �?             @       ������������������������       �                      @        ������������������������       �                      @        j       k                 ���E@ףp=
�?             $@       ������������������������       �                      @        l       m                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     :@        q                          @z6�>��?            y@       r       s                 ���@�o6�
�?�            �x@        ������������������������       �                     ;@        t                          @.�6�G,�?�             w@       u       �                    �?H?�߽��?�            �v@        v       �                    �?�\��N��?H            �\@        w       |                    �?,���i�?            �D@       x       {                 ���@      �?             @@        y       z                 0��@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     =@        }       ~                    @X�<ݚ�?             "@        ������������������������       �                      @               �                  S�2@և���X�?             @       �       �                    �?z�G�z�?             @        ������������������������       �                      @    o   �       �                 ���&@�q�q�?             @ ?��  ������������������������       �                     �?�]��  �       �                 �|Y=@      �?              @ [��  ������������������������       �                     �?a   y   ������������������������       �                     �?   
   ������������������������       �                      @e   t   �       �                    @:PZ(8?�?-            @R@    s   �       �                    @z�G�z�?             @ 6��  ������������������������       �                      @`W��  �       �                    @�q�q�?             @    d   ������������������������       �                     �?0 ��  ������������������������       �                      @   t   �       �                    ,@�t����?)             Q@    .   ������������������������       �                     $@       �       �                   �"@J�8���?$             M@    s   �       �                    @�ՙ/�?             5@Y��  �       �                    ;@���Q��?             4@(z�  �       �                    �?������?
             .@�z�  �       �                 pf� @d}h���?	             ,@��z�  �       �                   �7@�C��2(�?             &@ v��  ������������������������       �                     @����  �       �                 �&B@z�G�z�?             @ s�|�  ������������������������       �                     �?p��  ������������������������       �                     @p�I}�  �       �                    3@�q�q�?             @ ��  ������������������������       �                     �?p�a}�  ������������������������       �                      @����  ������������������������       �                     �?p7I}�  �       �                 �?� @z�G�z�?             @�2�  ������������������������       �                     @���  ������������������������       �                     �? �.}�  ������������������������       �                     �? &�|�  �       �                 03�1@��G���?            �B@���  �       �                    �?�X����?             6@J}�  �       �                     @ҳ�wY;�?             1@�2�  �       �                   �3@������?
             .@ g2�  ������������������������       �                     �?P���  �       �                   �0@d}h���?	             ,@�d}�  �       �                 �|�;@8�Z$���?             *@ H�z�  ������������������������       �                      @ .�|�  �       �                 ���.@���Q��?             @k��  �       �                    �?      �?             @�1�  �       �                   �@@      �?              @ ���  ������������������������       �                     �?��a}�  ������������������������       �                     �?���  ������������������������       �                      @Ps��  ������������������������       �                     �?Nz�  ������������������������       �                     �?�a}�  ������������������������       �                      @�a��  �       �                   �;@z�G�z�?             @ l��  ������������������������       �                     �?Е��  ������������������������       �                     @0 b}�  ������������������������       �                     .@�T��  �       �                 ��@H%u��?�            @o@ �z�  ������������������������       �                     @���  �       �                    #@0�v����?�            �n@ �z�  �       �                     @     ��?             0@ ���  ������������������������       �                     @����  �       �                    @ףp=
�?             $@��  �       �                    �?z�G�z�?             @ ��  ������������������������       �                     �?�:��  �       �                 ���A@      �?             @ c��  �       �                    @      �?              @ ���  ������������������������       �                     �?p�z�  ������������������������       �                     �? �z�  ������������������������       �                      @�<��  ������������������������       �                     @ x��  �       �                    �?,���>�?�            �l@ v,}�  �       �                 03�-@д>��C�?'             M@�'�  �       �                 �|Y=@ףp=
�?              I@ ��  �       �                   �<@�<ݚ�?             "@q��  ������������������������       �                     @�9��  ������������������������       �                      @ $b}�  �       �                 �|Y?@��p\�?            �D@V��  �       �                    �?ܷ��?��?             =@�4�  �       �                 ���@�����H�?             ;@ `��  ������������������������       �                     @P]��  �       �                 P�J@؇���X�?             5@c��  �       �                 ���@R���Q�?             4@ �G}�  �       �                    �?�����H�?             "@%b}�  ������������������������       �r�q��?             @��2�  ������������������������       �                     @ �z�  ������������������������       �"pc�
�?             &@ Q��  ������������������������       �                     �?���  ������������������������       �                      @p��  ������������������������       �                     (@0���  �       �                 ��.@      �?              @ �4�  ������������������������       �                     @�5��  �       �                    �?���Q��?             @ ���  ������������������������       �                     �?�z��  �       �                    �?      �?             @P��  ������������������������       �                     @@��  ������������������������       �                     �?����  �                         @@@���y�?p            �e@�z�  �                          �?D��*�4�?\            @a@j��  �                          �?�[|x��?U            �_@��  �       �                 �!&B@�H�@=��?M            �[@���  �       �                 �|�=@ �h�7W�?J            �Z@&b}�  �       �                 @3�@��8�$>�?C            @X@�4�  ������������������������       �        $             H@0v�|�  �       �                 @�!@Hm_!'1�?            �H@`��  �       �                   � @PN��T'�?             ;@�z�  �       �                 0S5 @�r����?             .@k��  �       �                   �3@؇���X�?             ,@ O�|�  �       �                    1@�q�q�?             @ v�|�  ������������������������       �                     �? v�|�  ������������������������       �                      @�b��  ������������������������       �                     &@h��  ������������������������       �                     �?h��  �       �                   �7@r�q��?             (@@��  ������������������������       �                      @0���  �       �                 �|Y<@      �?             @ s�|�  ������������������������       �                      @ s�|�  ������������������������       �                      @����  ������������������������       �                     6@ �z�  �       �                   �?@�<ݚ�?             "@�z�  �       �                   �>@���Q��?             @ ��  �       �                 �̌!@      �?              @ ��  ������������������������       �                     �?@��  ������������������������       �                     �?�e��  �       �                 pff@�q�q�?             @ ��|�  ������������������������       �                      @'�z�  ������������������������       �                     �?p���  ������������������������       �                     @ �4�  �       �                    ;@z�G�z�?             @ v��  ������������������������       �                      @p��|�                            >@�q�q�?             @ �z�  ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     .@        ������������������������       �                     (@        ������������������������       �                    �A@                               �:@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h*h-K ��h/��R�(KM	KK��h]�B�       �{@     �p@     �`@      f@      <@     �T@      .@      "@       @      "@       @      @              @       @                       @      *@              *@     �R@      "@     �Q@      @      N@      @      @              @      @      �?              �?      @               @     �J@             �B@       @      0@      �?      ,@      �?                      ,@      �?       @      �?                       @      @      &@      �?       @      �?                       @       @      @              @       @              @      @      @      �?              �?      @                       @     �Z@     �W@      @     �P@      �?      8@      �?                      8@       @      E@      �?      D@              8@      �?      0@      �?       @              �?      �?      �?      �?                      �?              ,@      �?       @      �?                       @     �Y@      <@     @S@      <@     @S@      7@     @P@      (@      ,@             �I@      (@     �D@      (@      =@      &@      &@      @      $@      @      $@      @      @      @      @      �?              �?      @                      @      @                      �?      �?              2@      @      0@      @      ,@      @       @      @       @       @      @       @               @      @              @                      �?      @               @      @      �?      �?      �?       @       @              (@      �?      @              @      �?      @                      �?      $@              (@      &@      @              @      &@      @       @       @               @       @               @       @              �?      "@               @      �?      �?      �?                      �?              @      :@             0s@     @W@     �r@     @W@      ;@             0q@     @W@      q@     �V@      K@      N@      @      B@      �?      ?@      �?       @               @      �?                      =@      @      @               @      @      @      @      �?       @               @      �?      �?              �?      �?              �?      �?                       @     �H@      8@      �?      @               @      �?       @      �?                       @      H@      4@      $@              C@      4@       @      *@       @      (@      @      &@      @      &@      �?      $@              @      �?      @      �?                      @       @      �?              �?       @              �?              @      �?      @                      �?              �?      >@      @      .@      @      &@      @      &@      @              �?      &@      @      &@       @       @              @       @      @      �?      �?      �?              �?      �?               @                      �?              �?               @      @      �?              �?      @              .@             �k@      >@              @     �k@      ;@      "@      @              @      "@      �?      @      �?      �?              @      �?      �?      �?      �?                      �?       @              @             `j@      4@      H@      $@     �F@      @      @       @      @                       @      C@      @      :@      @      8@      @      @              2@      @      1@      @       @      �?      @      �?      @              "@       @      �?               @              (@              @      @              @      @       @              �?      @      �?      @                      �?     `d@      $@      `@      $@      ]@      $@     @Y@      $@      Y@      @     @W@      @      H@             �F@      @      7@      @      *@       @      (@       @      �?       @      �?                       @      &@              �?              $@       @       @               @       @               @       @              6@              @       @      @       @      �?      �?      �?                      �?       @      �?       @                      �?      @              �?      @               @      �?       @      �?                       @      .@              (@             �A@              �?      @              @      �?              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�R�[hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B�C         \                    �?�s�ˈ.�?�           8�@      @       U                 p�H@�d�����?�            �l@              4                    �?Ҙ$�Ų�?k            �d@      @                            @�<ݚ�?=            �X@               
                    �?�(\����?             D@    �B@                          �J@�nkK�?             7@     ,@������������������������       �                     4@      &@       	                 `f�2@�q�q�?             @      @������������������������       �                     �?0i�y�  ������������������������       �                      @i�y�  ������������������������       �        
             1@i�y�                             �?:���W�?#            �M@ i�y�                             �?�+e�X�?             9@ i�y�                          H�%@���Q��?             $@ i�y�  ������������������������       �                     @ i�y�                          03�-@z�G�z�?             @ i�y�  ������������������������       �                     @      @                        �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?      @                        X�,A@�r����?             .@       ������������������������       �                     *@      @������������������������       �                      @      �?       /                    �?�ʻ����?             A@     �?       .                    �?*;L]n�?             >@     &@                           '@П[;U��?             =@       @������������������������       �                     @      �?                          �4@      �?             :@        ������������������������       �                     @     @W@       )                 `��!@\X��t�?             7@     ?@       (                    C@������?	             .@     =@        !                 P�@d}h���?             ,@      �?������������������������       �                     @      @"       '                 �|Y>@      �?              @       #       &                 �|�;@      �?             @     6@$       %                   �8@      �?              @      ,@������������������������       �                     �?      @������������������������       �                     �?      �?������������������������       �                      @        ������������������������       �                     @      @������������������������       �                     �?      �?*       +                    ;@      �?              @     >@������������������������       �                     @      �?,       -                   �@@�q�q�?             @        ������������������������       �                      @       @������������������������       �                     �?      @������������������������       �                     �?       @0       1                    @      �?             @      �?������������������������       �                     �?      �?2       3                 ��l4@�q�q�?             @      �?������������������������       �                     �?      @������������������������       �                      @      @5       <                     @�'�=z��?.            �P@      �?6       9                    6@؇���X�?             5@      �?7       8                 ��m1@      �?             @        ������������������������       �                      @        ������������������������       �                      @        :       ;                   �B@�IєX�?             1@     @������������������������       �                     0@      H@������������������������       �                     �?      @=       @                    �?f.i��n�?            �F@        >       ?                 ��.@�q�q�?             @        ������������������������       �                      @      �?������������������������       �                     @      7@A       J                 03�1@��Sݭg�?            �C@      &@B       I                    �?�q�q�?             (@     �?C       H                 ��Y.@���Q��?             $@       D       G                    �?z�G�z�?             @     6@E       F                    6@      �?             @      @������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        K       P                    @�>����?             ;@       L       O                 ���4@���7�?             6@        M       N                 03C3@�q�q�?             @       ������������������������       �                      @       ������������������������       �                     �?       ������������������������       �        
             3@       Q       R                 ��T?@z�G�z�?             @        ������������������������       �                      @        S       T                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        V       [                 ���Q@$Q�q�?+            �O@        W       X                    �?�J�4�?             9@       ������������������������       �                     3@        Y       Z                 ���P@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     C@        ]       �                    �?���A�
�?*           0~@        ^       k                 ��K.@N��c��?1            @S@        _       d                   �6@������?            �D@        `       a                    �?      �?             @        ������������������������       �                     �?        b       c                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        e       f                 �|=@�?�|�?            �B@        ������������������������       �                     &@        g       j                   @@ ��WV�?             :@       h       i                 ���@�C��2(�?             &@       ������������������������       �                     @        ������������������������       �      �?             @       ������������������������       �                     .@        l       w                    �?b�2�tk�?             B@       m       r                 �|Y<@�z�G��?             4@        n       q                    9@����X�?             @        o       p                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?       ������������������������       �                     @        s       v                   �F@$�q-�?
             *@        t       u                 X�,@@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @       x                           �?      �?             0@       y       |                 ��G@և���X�?
             ,@        z       {                 ��3@      �?              @        ������������������������       �                     @        ������������������������       �                     @        }       ~                 ���X@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?       ������������������������       �                      @        �       �                   �/@|g�&��?�            `y@       �       �                    �?<N_�U��?�            �p@���  �       �                 �?�@     �?�             p@ ���  �       �                     @������?M            �^@ z��  ������������������������       �                     &@    t   �       �                    �?�h����?E             \@    )   �       �                  ��@8�Z$���?             *@    e   ������������������������       �                      @   E   �       �                    �?"pc�
�?	             &@���  �       �                 �|Y=@�<ݚ�?             "@ v��  ������������������������       �                     �?    e   �       �                 ��(@      �?              @��  ������������������������       �r�q��?             @   e   ������������������������       �                      @       ������������������������       �                      @    '   �       �                   �7@��:x�ٳ?:            �X@    x   ������������������������       �                     A@����  �       �                 �Yu@����?&            @P@   "   �       �                 �&B@(N:!���?            �A@   j   �       �                   �8@`Jj��?             ?@    _   �       �                 �&b@���Q��?             @ S��  ������������������������       �                     @��  ������������������������       �                      @    s   ������������������������       �                     :@��  �       �                    �?      �?             @    p   ������������������������       �                      @ ���  ������������������������       �                      @   e   ������������������������       �                     >@���  �       �                   �0@���H��?N            �`@    _   �       �                 �̌!@�q�q�?             @    e   ������������������������       �                      @ ���  ������������������������       �                     �?   t   �       �                   �*@ ����?L            @`@   o   �       �                   �A@���5��?D            �\@8��  �       �                   �<@8�Z$���?7            �V@   m   �       �                   �3@$�q-�?             J@    t   �       �                     @������?	             .@    h   �       �                    &@      �?             @ {��  ������������������������       �      �?              @   o   ������������������������       �                      @e   x   �       �                   �1@���!pc�?             &@    e   ������������������������       �                     @\и�  �       �                 0S5 @և���X�?             @    t   ������������������������       �                     @@��  ������������������������       �                     @        ������������������������       �                    �B@`���  �       �                 ��)"@��Sݭg�?            �C@׸�  �       �                   �?@�KM�]�?             3@   n   �       �                   �>@8�Z$���?             *@       �       �                 �|Y=@�8��8��?
             (@ `��  ������������������������       �                     �?�и�  �       �                 ��) @�C��2(�?	             &@3��  ������������������������       �                     "@]   :   �       �                 pf� @      �?              @ ���  ������������������������       �                     �?   m   ������������������������       �                     �? ��  ������������������������       �                     �?    b   ������������������������       �                     @a��  �       �                 �|�=@���Q��?             4@ ���  ������������������������       �                     @       �       �                   �@@�t����?             1@���  �       �                    $@�θ�?	             *@ ���  �       �                   �?@      �?             @ b��  ������������������������       �                     @:��  ������������������������       �                     �?    u   ������������������������       �                     "@"   "   ������������������������       �      �?             @MU��  ������������������������       �                     7@�T��  ������������������������       �                     0@       �       �                    �?���|���?             &@   
   �       �                     @X�<ݚ�?             "@ Y��  ������������������������       �                     �? Ը�  �       �                   �*@      �?              @ ���  �       �                 xFT$@���Q��?             @        ������������������������       �                      @�t��  ������������������������       �                     @f   r   ������������������������       �                     @�ĸ�  ������������������������       �                      @ |��  �       �                    @4kMU*m�?X            `a@ Ǹ�  �       �                   �;@������?             .@        ������������������������       �                     @        �       �                    @      �?              @    p   ������������������������       �                     @       ������������������������       �                     @ o��  �                          �?���b��?P             _@��  �       �                    �? �&�T�?:             W@ո�  �       �                     @���3�E�?$             J@o��  �       �                 ��$:@�*/�8V�?             �G@        ������������������������       �        	             .@ ���  �       �                   �>@      �?             @@:��  �       �                 `fF<@�t����?             1@X��  �       �                    K@      �?             $@n��  �       �                 03k:@����X�?             @ ��  ������������������������       �                     �?���  �       �                 �|�<@�q�q�?             @    s   ������������������������       �                      @ i��  �       �                 X��B@      �?             @    -   ������������������������       �                     �?<���  �       �                   @G@�q�q�?             @   -   ������������������������       �      �?              @    -   ������������������������       �                     �?    -   ������������������������       �                     @�ĸ�  ������������������������       �                     @i   c   ������������������������       �                     .@ j��  �       �                 �|�>@���Q��?             @   -   �       �                 �T�C@�q�q�?             @    -   ������������������������       �                     �?   -   �       �                 �|�;@      �?              @ Ǹ�  ������������������������       �                     �?    m   ������������������������       �                     �?       ������������������������       �                      @ ���  �       �                    �?      �?             D@���  �       �                  x#J@r٣����?            �@@       ������������������������       �        
             1@   a   �       �                    F@      �?             0@��  �       �                 `f�K@�q�q�?             (@   l   �       �                    7@      �?              @        ������������������������       �                     @ ���  �       �                 `�iJ@z�G�z�?             @    n   ������������������������       �                      @ ���  �       �                    @@�q�q�?             @ e��  ������������������������       �                      @   _   ������������������������       �                     �?   g   ������������������������       �                     @ ��  ������������������������       �                     @   r   �       �                 �|�:@����X�?             @ R��  ������������������������       �                     @   r                               @�q�q�?             @    p   ������������������������       �                     �?        ������������������������       �                      @                                 @      �?             @@                                �?`Jj��?             ?@                                 @�X�<ݺ?             2@        ������������������������       �                     @              
                   @@4և���?	             ,@             	                   0@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                 �?$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     �?        �t�bh�h*h-K ��h/��R�(KMKK��h]�B�       �|@     @o@      N@      e@      L@     @[@      6@     @S@      �?     �C@      �?      6@              4@      �?       @      �?                       @              1@      5@      C@      @      3@      @      @              @      @      �?      @              �?      �?              �?      �?               @      *@              *@       @              .@      3@      *@      1@      *@      0@              @      *@      *@      @              $@      *@      @      &@      @      &@              @      @      @      @      �?      �?      �?      �?                      �?       @                      @      �?              @       @      @              �?       @               @      �?                      �?       @       @              �?       @      �?              �?       @              A@      @@      @      2@       @       @               @       @              �?      0@              0@      �?              ?@      ,@       @      @       @                      @      =@      $@      @       @      @      @      @      �?      @      �?              �?      @              �?                      @               @      9@       @      5@      �?       @      �?       @                      �?      3@              @      �?       @               @      �?              �?       @              @     �M@      @      5@              3@      @       @               @      @                      C@     y@     �T@     �M@      2@     �B@      @      �?      @              �?      �?       @               @      �?              B@      �?      &@              9@      �?      $@      �?      @              @      �?      .@              6@      ,@      ,@      @       @      @       @      �?       @                      �?              @      (@      �?      @      �?      @                      �?       @               @       @      @       @      @      @              @      @              �?      @              @      �?               @             `u@      P@      n@      :@     @m@      6@     @]@      @      &@             �Z@      @      &@       @       @              "@       @      @       @              �?      @      �?      @      �?       @               @             �W@      @      A@             �N@      @      ?@      @      =@       @      @       @      @                       @      :@               @       @               @       @              >@             @]@      0@      �?       @               @      �?              ]@      ,@      Y@      ,@     @S@      ,@      H@      @      &@      @      @      �?      �?      �?       @               @      @      @              @      @              @      @             �B@              =@      $@      1@       @      &@       @      &@      �?      �?              $@      �?      "@              �?      �?              �?      �?                      �?      @              (@       @              @      (@      @      $@      @      �?      @              @      �?              "@               @       @      7@              0@              @      @      @      @              �?      @      @       @      @       @                      @      @               @             @Y@      C@      @      &@              @      @      @              @      @             @X@      ;@     �P@      9@     �B@      .@     �A@      (@      .@              4@      (@      @      (@      @      @       @      @              �?       @      @               @       @       @      �?              �?       @      �?      �?              �?      @                      @      .@               @      @       @      �?      �?              �?      �?              �?      �?                       @      >@      $@      9@       @      1@               @       @      @       @      @      @      @              �?      @               @      �?       @               @      �?                      @      @              @       @      @              �?       @      �?                       @      >@       @      =@       @      1@      �?      @              *@      �?       @      �?              �?       @              @              (@      �?              �?      (@              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�v}hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtK�huh*h-K ��h/��R�(KK���h|�B@?         b                    �?��eC~�?�           8�@     @S@       ]                 p�H@������?�            `n@              D                    �?�H�]�r�?p            @e@���         	                 ��@r�0p�?F            �Z@                                   �?P���Q�?             4@       ������������������������       �        	             ,@      3@                        ���@r�q��?             @     *@������������������������       �                     @      &@������������������������       �                     �?        
                            @��V#�?8            �U@                                   L@>A�F<�?             C@     4@                           �?     ��?             @@      @������������������������       �                     @      ,@                        `f�)@�����H�?             ;@        ������������������������       �                     &@      �?                           �?     ��?             0@     �?                           :@r�q��?             (@      @������������������������       �                      @        ������������������������       �                     $@                                   <@      �?             @      @                          �9@      �?              @        ������������������������       �                     �?      @������������������������       �                     �?      �?������������������������       �                      @     �?                        `f�2@�q�q�?             @      &@������������������������       �                     @       @������������������������       �                      @      �?       7                 �|�<@     ��?              H@              ,                 Ь�!@�5��?             ;@    @W@       #                   �6@���Q��?             .@      ?@       "                 �&B@�<ݚ�?             "@      =@        !                    4@      �?             @      �?������������������������       �                      @      @������������������������       �                      @        ������������������������       �                     @      �?$       %                 �&B@�q�q�?             @      @������������������������       �                     �?       @&       '                   �9@���Q��?             @        ������������������������       �                      @        (       )                   �@�q�q�?             @        ������������������������       �                     �?      @*       +                 �?�@      �?              @        ������������������������       �                     �?      @������������������������       �                     �?       @-       0                    �?r�q��?	             (@      �?.       /                    4@�q�q�?             @        ������������������������       �                     �?      @������������������������       �                      @      @1       6                 ��.@�����H�?             "@       2       3                   �-@z�G�z�?             @      �?������������������������       �                      @      @4       5                 �yG(@�q�q�?             @     &@������������������������       �                      @        ������������������������       �                     �?      (@������������������������       �                     @      @8       =                 �|Y>@���N8�?             5@      @9       :                    �?@4և���?             ,@     �?������������������������       �                     $@        ;       <                    �?      �?             @      �?������������������������       �                     �?      $@������������������������       �                     @       @>       A                    @@և���X�?             @       @?       @                    �?      �?             @      @������������������������       �                     �?       @������������������������       �                     @      @B       C                   �A@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        E       J                    �?      �?*             P@        F       I                    �?���Q��?	             .@       G       H                 `�@1@�eP*L��?             &@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        K       L                    @Rg��J��?!            �H@        ������������������������       �                     @        M       N                    (@��6���?             E@        ������������������������       �                      @        O       P                   �:@�ʻ����?             A@        ������������������������       �        
             &@        Q       \                     @�LQ�1	�?             7@       R       [                    @X�<ݚ�?
             2@       S       T                   �?@��.k���?	             1@        ������������������������       �                     @        U       V                     @�q�q�?             (@        ������������������������       �                     @        W       X                    �?      �?              @        ������������������������       �                      @        Y       Z                 ��p@@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ^       _                    !@��pBI�?0            @R@        ������������������������       �                     �?        `       a                    @�k~X��?/             R@       ������������������������       �        .            �Q@        ������������������������       �                     �?        c       n                    @K�(i�?"           @}@        d       i                    �?8����?             7@       e       f                     @�q�q�?             (@       ������������������������       �                     @        g       h                 �y�-@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        j       k                     @"pc�
�?             &@       ������������������������       �                     @        l       m                 pf�@@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        o       �                    �?4�<����?           �{@        p       {                 P�J.@����X�?4             U@        q       r                   @@     ��?             @@       ������������������������       �                     1@        s       z                 �(@z�G�z�?             .@        t       y                 �y�#@և���X�?             @       u       x                 �� @z�G�z�?             @       v       w                    ?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        |       �                    �?�E��
��?              J@       }       �                   �H@j���� �?            �I@       ~       �                     @      �?             E@              �                     �?��%��?            �B@       �       �                   �8@*;L]n�?             >@        �       �                  D�U@r�q��?             @    o   ������������������������       �                     �? ?��  ������������������������       �                     @�]��  �       �                    �?�q�q�?             8@[��  �       �                 �ܵ<@      �?             4@    y   ������������������������       �                      @   
   �       �                    �?r�q��?
             2@   t   �       �                 `f�A@      �?             (@    s   ������������������������       �                     @ 6��  �       �                 @�6M@      �?             @ W��  ������������������������       �                     @    d   ������������������������       �                     @0 ��  ������������������������       �                     @   t   �       �                 @��v@      �?             @   .   ������������������������       �                     @       ������������������������       �                     �?    s   ������������������������       �                     @Y��  �       �                    �?z�G�z�?             @ (z�  ������������������������       �                     �?�z�  ������������������������       �                     @��z�  ������������������������       �                     "@ v��  ������������������������       �                     �?����  �       �                 `ff:@���5���?�            �v@s�|�  �       �                    �?��S�jC�?�            pr@��  �       �                    )@(�s���?�            �o@ �I}�  ������������������������       �                      @ ��  �       �                   @E@ ��GS=�?�            @o@�a}�  �       �                   �D@�IєX�?�            �k@���  �       �                 ���@�X�<ݺ?�             k@ 7I}�  ������������������������       �                    �C@�2�  �       �                 �?$@ ,��-�?i             f@ ���  �       �                   �;@�㙢�c�?             7@ �.}�  ������������������������       �                     @ &�|�  �       �                    �?������?
             1@���  �       �                 �|Y=@d}h���?             ,@ J}�  ������������������������       �                      @�2�  ������������������������       ��8��8��?             (@ g2�  �       �                 �|Y?@�q�q�?             @ ���  ������������������������       �                     �?�d}�  ������������������������       �                      @ H�z�  �       �                 �?�@�kb97�?[            @c@ .�|�  ������������������������       �                    �A@k��  �       �                   �3@T(y2��?C            �]@ �1�  �       �                   �1@��2(&�?             6@ ���  ������������������������       �                     @��a}�  �       �                 0S5 @z�G�z�?	             .@ ��  �       �                   �2@      �?             @ s��  ������������������������       �                     �?Nz�  ������������������������       ��q�q�?             @�a}�  ������������������������       �                     &@�a��  �       �                    �?h�a��?7            @X@l��  �       �                 �|�=@ rpa�?5            @W@���  �       �                 @3�!@��v$���?!            �N@  b}�  �       �                 pf� @�nkK�?             7@T��  ������������������������       �        
             4@ �z�  �       �                    8@�q�q�?             @ ���  ������������������������       �                      @ �z�  ������������������������       �                     �? ���  ������������������������       �                     C@����  �       �                   �?@      �?             @@ ��  �       �                     @�<ݚ�?             "@ ��  ������������������������       �                     @�:��  �       �                 @3�@      �?             @ c��  ������������������������       �                     �? ���  �       �                 �̌!@�q�q�?             @ �z�  ������������������������       �                      @ �z�  ������������������������       �                     �?�<��  �       �                   �@@���}<S�?             7@ x��  ������������������������       �                     "@ v,}�  �       �                     @؇���X�?	             ,@�'�  �       �                   �3@؇���X�?             @��  �       �                   �A@r�q��?             @ q��  ������������������������       ��q�q�?             @�9��  ������������������������       �                     @ $b}�  ������������������������       �                     �?V��  �       �                 @3�@؇���X�?             @ �4�  ������������������������       ��q�q�?             @ `��  ������������������������       �                     @P]��  ������������������������       �                     @c��  �       �                 ���%@z�G�z�?             @ �G}�  ������������������������       �                     @%b}�  ������������������������       �      �?              @��2�  ������������������������       �                     =@ �z�  �       �                     @ qP��B�?            �E@ Q��  ������������������������       �                      @���  �       �                   �/@��?^�k�?            �A@��  ������������������������       �                     2@0���  �       �                    )@�IєX�?             1@ �4�  ������������������������       �                     �?�5��  ������������������������       �        
             0@ ���  �       �                    �?:ɨ��?-            �P@z��  �       �                    �?���Q��?              I@P��  �       �                     �?��.k���?             A@��  �       �                   �>@X�<ݚ�?             ;@���  �       �                    R@����X�?             5@�z�  �       �                   @=@�q�q�?             2@j��  �       �                 �|�<@���Q��?             $@ ��  ������������������������       �                     �?���  �       �                 `f�;@�q�q�?             "@&b}�  �       �                 �|�?@      �?              @ �4�  ������������������������       �                     @0v�|�  �       �                   �J@���Q��?             @ `��  ������������������������       �                     @�z�  ������������������������       �                      @k��  ������������������������       �                     �? O�|�  ������������������������       �                      @ v�|�  ������������������������       �                     @ v�|�  ������������������������       �                     @�b��  �       �                 �|�>@؇���X�?             @��  ������������������������       �                     @h��  ������������������������       �                     �?@��  �       �                 ��9L@      �?
             0@���  �       �                   �C@ףp=
�?             $@ s�|�  ������������������������       �                     @ s�|�  �       �                    G@�q�q�?             @���  �       �                     �?      �?              @ �z�  ������������������������       �                     �?�z�  ������������������������       �                     �? ��  ������������������������       �                     �? ��  �       �                   �D@      �?             @��  �       �                     �?      �?             @e��  ������������������������       �                     @ ��|�  ������������������������       �                     �?'�z�  ������������������������       �                      @p���  ������������������������       �                     0@ �4�  �t�b��     h�h*h-K ��h/��R�(KK�KK��h]�B�       p|@      p@     �O@     �f@     �N@     @[@      =@     @S@      �?      3@              ,@      �?      @              @      �?              <@      M@      @      ?@      @      =@              @      @      8@              &@      @      *@       @      $@       @                      $@      �?      @      �?      �?              �?      �?                       @      @       @      @                       @      5@      ;@      0@      &@      @      "@       @      @       @       @       @                       @              @      @       @      �?              @       @       @              �?       @              �?      �?      �?      �?                      �?      $@       @       @      �?              �?       @               @      �?      @      �?       @               @      �?       @                      �?      @              @      0@      �?      *@              $@      �?      @      �?                      @      @      @      @      �?              �?      @              �?       @               @      �?              @@      @@      "@      @      @      @      @                      @      @              7@      :@              @      7@      3@       @              .@      3@              &@      .@       @      $@       @      "@       @      @              @       @              @      @      @       @               @      @              @       @              �?              @               @     �Q@      �?              �?     �Q@             �Q@      �?             �x@      S@      @      0@      @      @              @      @       @               @      @               @      "@              @       @      @              @       @             x@      N@      N@      8@      =@      @      1@              (@      @      @      @      @      �?       @      �?              �?       @               @                       @       @              ?@      5@      >@      5@      5@      5@      4@      1@      *@      1@      @      �?              �?      @               @      0@      @      .@       @              @      .@      @      "@              @      @      @      @                      @              @      @      �?      @                      �?      @              �?      @      �?                      @      "@              �?             Pt@      B@     pq@      0@     �m@      .@               @     �m@      *@      j@      *@     �i@      (@     �C@             �d@      (@      3@      @      @              *@      @      &@      @               @      &@      �?       @      �?              �?       @             @b@       @     �A@             �[@       @      3@      @      @              (@      @      �?      @              �?      �?       @      &@              W@      @      V@      @      N@      �?      6@      �?      4@               @      �?       @                      �?      C@              <@      @      @       @      @               @       @              �?       @      �?       @                      �?      5@       @      "@              (@       @      @      �?      @      �?       @      �?      @              �?              @      �?       @      �?      @              @              @      �?      @              �?      �?      =@              E@      �?       @              A@      �?      2@              0@      �?              �?      0@              G@      4@      >@      4@      2@      0@      (@      .@      @      .@      @      (@      @      @              �?      @      @      @      @      @               @      @              @       @              �?                       @              @      @              @      �?      @                      �?      (@      @      "@      �?      @               @      �?      �?      �?              �?      �?              �?              @      @      �?      @              @      �?               @              0@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJg}�XhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMChuh*h-K ��h/��R�(KMC��h|�B�P         r                 `f�$@��t���?�           8�@      @                            @z�G�z�?�            @p@  o u r ������������������������       �                      @      =@       k                   @@@Z���c��?�            �o@     *@                            �?�۲I <�?�            �j@      @                        �|Y=@T�7�s��?#            �L@       @                        ���@"pc�
�?             &@      ;@       	                   �2@�q�q�?             @       @������������������������       �                     �?       
                        �{@      �?              @        ������������������������       �                     �?       ������������������������       �                     �?       ������������������������       �                      @                                03@�LQ�1	�?             G@                               ���@���"͏�?            �B@                                   �?$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@                                   �?�q�q�?             8@     @                        ��@�LQ�1	�?             7@      &@������������������������       �                      @                                   �?����X�?             5@                                  �?�q�q�?             2@        ������������������������       �                     @     �Q@                        ���@؇���X�?	             ,@      0@������������������������       �                     �?       @������������������������       �8�Z$���?             *@      @������������������������       �                     @      8@������������������������       �                     �?      @                           �?�<ݚ�?             "@       ������������������������       �                     @      5@������������������������       �                      @      1@!       4                    �?�IA��?e            �c@        "       3                 �|Y>@     ��?             0@       #       2                    �?���Q��?             .@       $       -                   �6@և���X�?             ,@       %       ,                 xF� @X�<ݚ�?             "@       &       +                    �?r�q��?             @       '       *                   �3@z�G�z�?             @        (       )                 P��@      �?              @        ������������������������       �                     �?       ������������������������       �                     �?       ������������������������       �                     @       ������������������������       �                     �?       ������������������������       �                     @       .       /                 �&B@z�G�z�?             @        ������������������������       �                      @       0       1                    9@�q�q�?             @       ������������������������       �                      @       ������������������������       �                     �?       ������������������������       �                     �?       ������������������������       �                     �?       5       H                 �?�@`	�<��?V            �a@       6       E                   �?@��p\�?.            �T@       7       <                 ���@ �\���?,            �S@        8       9                    7@����X�?             @        ������������������������       �                     @       :       ;                 �&b@      �?             @       ������������������������       �                      @       ������������������������       �                      @       =       D                 �?$@������?'             R@        >       ?                 �|Y;@HP�s��?             9@       ������������������������       �        
             2@        @       C                 �|Y>@����X�?             @       A       B                 ��@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                    �G@        F       G                   �@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        I       R                 @3�@��$�4��?(            �M@        J       Q                    �?X�<ݚ�?             "@       K       P                    �?      �?              @       L       M                   �9@և���X�?             @        ������������������������       �                      @        N       O                   �?@���Q��?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     �?        S       h                 �|�=@j�q����?"             I@       T       a                 @�!@��0{9�?             �G@       U       ^                   � @"pc�
�?            �@@       V       ]                 0S5 @�>4և��?             <@       W       \                   �4@�+$�jP�?             ;@        X       Y                    1@X�<ݚ�?             "@        ������������������������       �      �?             @        Z       [                   �2@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     2@        ������������������������       �                     �?        _       `                   �7@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        b       c                 ���"@@4և���?
             ,@        ������������������������       �                     @        d       e                   �<@ףp=
�?             $@       ������������������������       �                     @        f       g                 �|Y=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        i       j                    ?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        l       m                   @C@P�Lt�<�?             C@        ������������������������       �                     3@        n       o                    �?�}�+r��?             3@        ������������������������       �                      @        p       q                   �C@�IєX�?
             1@        ������������������������       ��q�q�?             @        ������������������������       �                     ,@        s                           @.iI\��?           0|@       t       �                  x#J@$;hB��?�            @s@       u       �                   �<@��U��?�            �j@        v       �                    �?��V#�?1            �U@       w       x                    �?@3����?             K@        ������������������������       �                      @        y       �                    �?��<b�ƥ?             G@        z       {                   �6@�nkK�?	             7@        ������������������������       �                     "@        |                          �9@@4և���?             ,@        }       ~                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     7@    )   �       �                    �?     ��?             @@ D]i 
 ��       �                    �?և���X�?             @   .   �       �                   �8@���Q��?             @   t   �       �                 hf:@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?   g   ������������������������       �                      @    "   ������������������������       �                      @       �       �                   �>@HP�s��?             9@   f   ������������������������       �                     7@.   s   ������������������������       �                      @   b   �       �                    �?b����?R            �_@       �       �                  �?@�8�Վ��?Q            @_@       �       �                    �?D��ٝ�?B            @Y@        �       �                    �?�eP*L��?             6@    b   �       �                    D@r�q��?             @   _   ������������������������       �                     @        ������������������������       �                     �?       �       �                   @C@     ��?	             0@   t   �       �                 ��";@r�q��?             (@       �       �                   @@@�q�q�?             @    =   ������������������������       �                     @   p   �       �                   �A@�q�q�?             @    
   ������������������������       �                      @    s   ������������������������       �                     �?    =   ������������������������       �                     @       �       �                     �?      �?             @    s   ������������������������       �                     @    u   ������������������������       �                     �?        �       �                    �?���%&�?5            �S@   e   �       �                   �F@^H���+�?2            �R@   s   �       �                   @F@�[�IJ�?             �G@   e   �       �                   @E@�lg����?            �E@       �       �                     �?�e����?            �C@    r   �       �                 �|�?@�q�q�?             @   n   �       �                   �>@z�G�z�?             @   s   �       �                 `f�;@      �?              @        ������������������������       �                     �?o   k   ������������������������       �                     �?       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �C@4���C�?            �@@   e   �       �                   @B@����"�?             =@   n   �       �                    �?
;&����?             7@    o   ������������������������       �                     "@        �       �                    1@؇���X�?             ,@       �       �                   �'@�<ݚ�?             "@    l   ������������������������       �                     @   b   �       �                    @@�q�q�?             @    o   ������������������������       �                     @       ������������������������       ��q�q�?             @   h   ������������������������       �                     @    g   ������������������������       �                     @   w   �       �                   �,@      �?             @        ������������������������       �      �?              @    e   ������������������������       �                      @    N   ������������������������       �                     @o   n   ������������������������       �                     @    t   �       �                   �R@�<ݚ�?             ;@   H   �       �                    �?���B���?             :@    ,   ������������������������       �                     @    a   �       �                    �?���}<S�?             7@       �       �                   �I@�C��2(�?             6@   e   �       �                 ��:@r�q��?             (@       ������������������������       �                      @    r   �       �                 `f�;@      �?             @   P   ������������������������       �                      @        ������������������������       �                      @    k   ������������������������       �                     $@   e   ������������������������       �                     �?   e   ������������������������       �                     �?    a   �       �                    �?z�G�z�?             @    c   ������������������������       �                     �?    e   ������������������������       �                     @    a   �       �                    �?      �?             8@        ������������������������       �                     @l   a   ������������������������       �                     5@    n   ������������������������       �                     �?    v   �                         �O@�q�q�?A             X@   a   �       �                   �5@���!pc�?>             V@    c   �       �                   �1@��.k���?             1@   s   �       �                 ��f`@؇���X�?             @   i   ������������������������       �                     @    e   �       �                    �?      �?              @    x   ������������������������       �                     �?       ������������������������       �                     �?   n   �       �                    �?z�G�z�?             $@   l   ������������������������       �                      @        ������������������������       �                      @   a   �       �                 `fmj@@���?T�?3            �Q@       �       �                    �?     8�?.             P@       �       �                 ���P@���-T��?-             O@    h   �       �                 03sP@�z�G��?             4@   a   �       �                    �?@�0�!��?             1@        ������������������������       �                     $@   e   �       �                   �H@և���X�?             @       �       �                    �?z�G�z�?             @    I   ������������������������       �                     @       �       �                 0�nL@      �?              @        ������������������������       �                     �?   c   ������������������������       �                     �?    a   ������������������������       �                      @    f   ������������������������       �                     @        �       �                    �?@4և���?              E@   e   �       �                    �?@-�_ .�?            �B@   o   �       �                    �?`Jj��?             ?@   "   ������������������������       �                     0@    o   �       �                    �?�r����?             .@    ,   ������������������������       �                     @       �       �                   �H@      �?              @   e   �       �                 ЈT@؇���X�?             @    E   ������������������������       �                     @    _   �       �                   �D@      �?             @    e   ������������������������       �                      @   x   �       �                 Ј�U@      �?              @    ,   ������������������������       �                     �?    h   ������������������������       �                     �?    
   ������������������������       �                     �?        ������������������������       �                     @   o   �       �                 ��W@z�G�z�?             @    t   ������������������������       �                     @    t   ������������������������       �                     �?"   
   ������������������������       �                      @    t   �       �                    �?և���X�?             @        ������������������������       �                     �?    ,   �                          �?      �?             @   s                          �̾w@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @                                 �?x�f��^�?[            �a@                                 �?�>$�*��?            �D@                             X�,A@��+7��?             7@             	                  �0@��s����?             5@        ������������������������       �                     @        
                        �7@������?             .@        ������������������������       �                     �?                              �|Y=@d}h���?             ,@        ������������������������       �                      @                                 �?      �?             (@                              S�-@�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @                                 �?�q�q�?             2@                             03�-@�eP*L��?             &@                                 3@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                                 �?r�q��?             @                                �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @              8                   �?t�F�}�?B            �Y@              /                   �?�q�q�?'             N@        !      *                ���5@*;L]n�?             >@       "      )                  �D@     ��?
             0@       #      (                   7@�r����?	             .@        $      '                   �?      �?             @       %      &                   +@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     �?        +      .                  @C@����X�?             ,@        ,      -                X��@@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        0      1                   )@������?             >@        ������������������������       �                     @        2      7                   ;@H%u��?             9@        3      6                   �?և���X�?             @        4      5                �!&B@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     2@        9      B                   @@4և���?             E@        :      ;                   �?���!pc�?             &@        ������������������������       �                     @        <      =                   @և���X�?             @        ������������������������       �                     @        >      ?                   �?      �?             @        ������������������������       �                      @        @      A                ��T?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ?@        �t�bh�h*h-K ��h/��R�(KMCKK��h]�B0       �{@     �p@      j@      J@       @              i@      J@     `d@     �I@      @@      9@       @      "@       @      �?      �?              �?      �?      �?                      �?               @      >@      0@      <@      "@      (@      �?              �?      (@              0@       @      .@       @               @      .@      @      (@      @              @      (@       @      �?              &@       @      @              �?               @      @              @       @             ``@      :@      "@      @      "@      @       @      @      @      @      �?      @      �?      @      �?      �?              �?      �?                      @              �?      @              @      �?       @               @      �?       @                      �?      �?                      �?     �^@      3@      S@      @     �R@      @      @       @      @               @       @       @                       @     �Q@       @      7@       @      2@              @       @      @       @      @                       @       @             �G@              �?       @               @      �?              G@      *@      @      @      @      @      @      @       @               @      @              �?       @       @              �?      �?             �D@      "@      D@      @      ;@      @      7@      @      6@      @      @      @      @      �?      �?      @               @      �?       @      2@              �?              @      �?      @                      �?      *@      �?      @              "@      �?      @               @      �?              �?       @              �?       @               @      �?             �B@      �?      3@              2@      �?       @              0@      �?       @      �?      ,@             @m@      k@     �a@     �d@     �[@     �Y@      <@      M@      �?     �J@               @      �?     �F@      �?      6@              "@      �?      *@      �?      @      �?                      @              "@              7@      ;@      @      @      @       @      @       @      �?       @                      �?               @       @              7@       @      7@                       @     �T@      F@     �T@     �E@     �N@      D@      (@      $@      �?      @              @      �?              &@      @      $@       @      @       @      @              �?       @               @      �?              @              �?      @              @      �?             �H@      >@      H@      :@      ;@      4@      ;@      0@      7@      0@      @       @      @      �?      �?      �?      �?                      �?      @                      �?      3@      ,@      2@      &@      (@      &@              "@      (@       @      @       @      @              @       @      @              �?       @      @              @              �?      @      �?      �?               @      @                      @      5@      @      5@      @              @      5@       @      4@       @      $@       @       @               @       @               @       @              $@              �?                      �?      �?      @      �?                      @      5@      @              @      5@                      �?      @@      P@      8@      P@      "@       @      �?      @              @      �?      �?      �?                      �?       @       @       @                       @      .@      L@      &@     �J@      "@     �J@      @      ,@      @      ,@              $@      @      @      �?      @              @      �?      �?              �?      �?               @              @              @     �C@       @     �A@       @      =@              0@       @      *@              @       @      @      �?      @              @      �?      @               @      �?      �?      �?                      �?      �?                      @      �?      @              @      �?               @              @      @      �?              @      @      @       @      @                       @              �?       @              W@     �I@      2@      7@      @      1@      @      1@              @      @      &@      �?              @      &@               @      @      "@      @      @      @                      @               @       @              (@      @      @      @      @      �?              �?      @              �?      @      �?      �?      �?                      �?              @      @             �R@      <@     �A@      9@      *@      1@      @      *@       @      *@       @       @       @      �?              �?       @                      �?              &@      �?              $@      @      @      @      @                      @      @              6@       @              @      6@      @      @      @      �?      @      �?                      @      @              2@             �C@      @       @      @      @              @      @      @              �?      @               @      �?      �?      �?                      �?      ?@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ	�tlhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B@D         J                    �?�4�O��?�           8�@               5                    �?r�=���?~            �h@                                  �?T �����?[             c@       @                           �?�i�y�?$            �O@    �M@                           �?`Ӹ����?            �F@       @������������������������       �                     6@      @                            @���}<S�?             7@        ������������������������       �                     @        	       
                 ���@�����H�?             2@ T��  ������������������������       �                      @pO��  ������������������������       �        
             0@�_��  ������������������������       �        
             2@�W��                              �?��Hg���?7            �V@ _��                             �?և���X�?             5@]��                             �?���Q��?             4@���                          `f�A@�q�q�?             (@P��  ������������������������       �                     @      �?������������������������       �                     @                                  �5@      �?              @      �?������������������������       �                      @                                  �H@r�q��?             @     �?������������������������       �                     @      3@������������������������       �                     �?      C@������������������������       �                     �?      @                        ���@�~t��?*            @Q@        ������������������������       �        
             2@      �?       4                    �?��x_F-�?             �I@     ,@       3                 �|�=@j�q����?             I@              *                    �?      �?             B@     �?       %                   �:@���y4F�?             3@       @                         �&�)@�q�q�?             @        ������������������������       �                     �?        !       "                   �8@z�G�z�?             @ ���  ������������������������       �                     @�8��  #       $                 �0@      �?              @ ���  ������������������������       �                     �?0���  ������������������������       �                     �?���  &       )                   @@8�Z$���?             *@ >��  '       (                 �|=@�q�q�?             @ ��  ������������������������       �                      @p��  ������������������������       �      �?             @0��  ������������������������       �                     @��  +       .                 �|Y=@�t����?
             1@ ��  ,       -                  ��@      �?             @ ���  ������������������������       �                      @     �?������������������������       �                      @���  /       2                    �?�θ�?             *@��  0       1                  s�@�z�G��?             $@ ���  ������������������������       �                     @(N��  ������������������������       �      �?             @0���  ������������������������       �                     @      @������������������������       �                     ,@ ���  ������������������������       �                     �?���  6       C                    �?8�A�0��?#             F@���  7       <                 �|Y=@�LQ�1	�?             7@���  8       ;                 03�-@r�q��?
             (@ ��  9       :                    &@�q�q�?             @ ���  ������������������������       �                     �? ���  ������������������������       �                      @0��  ������������������������       �                     "@0<��  =       B                    �?�eP*L��?	             &@���  >       ?                   @E@r�q��?             @ ���  ������������������������       �                     @b��  @       A                 <3gH@�q�q�?             @ ��  ������������������������       �                     �?       @������������������������       �                      @      �?������������������������       �                     @      �?D       I                     @؇���X�?             5@       E       H                 �̾w@�θ�?             *@       F       G                    )@�C��2(�?
             &@        ������������������������       �                     �?        ������������������������       �        	             $@        ������������������������       �                      @        ������������������������       �                      @        K       �                    �?D����?C           �@        L       m                    �?�BA����?f            `d@        M       l                   �J@�7�QJW�?/            �R@       N       [                     @v���a�?.            @R@       O       P                   �6@$�q-�?             J@        ������������������������       �        	             2@        Q       Z                   �*@�t����?             A@        R       S                   �'@�	j*D�?
             *@        ������������������������       �                      @        T       U                    :@���|���?             &@        ������������������������       �                      @        V       W                   �B@�<ݚ�?             "@       ������������������������       �                     @        X       Y                    D@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     5@        \       k                    @�q�q�?             5@       ]       j                 @�"@�z�G��?             4@       ^       i                 `��!@և���X�?
             ,@       _       b                 ���@�q�q�?	             (@        `       a                 �|Y:@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        c       d                    4@և���X�?             @        ������������������������       �                      @        e       f                 @3�@z�G�z�?             @       ������������������������       �                     @        g       h                 �|Y>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        n       �                 �D�H@��7��?7             V@       o       �                    @�{r٣��?'            �P@       p       q                    @JJ����?            �G@        ������������������������       �                     @        r       �                    �?�D����?             E@       s       �                    @\�Uo��?             C@       t       u                   �6@և���X�?            �A@        ������������������������       �                     @        v       }                     @     ��?             @@        w       x                   �7@      �?             (@        ������������������������       �                      @        y       |                    �?ףp=
�?             $@       z       {                    D@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ~                        �|Y=@�z�G��?             4@        ������������������������       �                     @        �       �                    �?���Q��?             .@        �       �                 ��1@�q�q�?             @       ������������������������       �                     @    p   ������������������������       �                      @    s   �       �                 `fV6@�<ݚ�?             "@    f   ������������������������       �                     �?        �       �                 ��T?@      �?              @       ������������������������       �                     @        ������������������������       �                     �?    n   ������������������������       �                     @        �       �                    �?      �?             @    o   ������������������������       �                      @    t   ������������������������       �                      @        �       �                 pfv2@p�ݯ��?
             3@        ������������������������       �                     @   s   �       �                    �?$�q-�?             *@    S   ������������������������       �                      @       �       �                 ��T?@z�G�z�?             @   T   ������������������������       �                     @   t   ������������������������       �                     �?   y   �       �                    #@�C��2(�?             6@    t   ������������������������       �                     �?        �       �                 ���P@���N8�?             5@    ,   ������������������������       �                     $@    y   �       �                 X�,@@�C��2(�?             &@        �       �                    �?�q�q�?             @    o   ������������������������       �                     �?       �       �                 ���d@      �?              @    n   ������������������������       �                     �?   m   ������������������������       �                     �?    i   ������������������������       �                      @        �       �                     �?PN��T'�?�            �u@    e   �       �                   �>@�j�'�=�?*            �P@    
   �       �                   �<@r�q��?             8@        ������������������������       �                     @   _   �       �                   �Q@��Q��?             4@       �       �                   @E@�E��ӭ�?             2@       �       �                 03:@d}h���?
             ,@    i   ������������������������       �                      @    y   �       �                 03k:@      �?             @        ������������������������       �                     �?    n   �       �                 �|�?@���Q��?             @   o   �       �                 `fF<@      �?             @    b   ������������������������       �                      @       �       �                 �|Y=@      �?              @        ������������������������       �                     �?   t   ������������������������       �                     �?       ������������������������       �                     �?       �       �                    K@      �?             @   l   �       �                   @G@�q�q�?             @   .   ������������������������       �      �?              @    n   ������������������������       �                     �?       ������������������������       �                     �?        ������������������������       �                      @        �       �                 �|�<@��s����?             E@        ������������������������       �                     @    v   �       �                    �?�ݜ�?            �C@       �       �                   �E@4?,R��?             B@       �       �                  x#J@�E��ӭ�?             2@       ������������������������       �                     "@    e   �       �                 �|Y>@X�<ݚ�?             "@    a   ������������������������       �                      @        �       �                 `f�K@����X�?             @    v   �       �                 `�iJ@�q�q�?             @        ������������������������       �                     �?       ������������������������       �                      @   F   ������������������������       �                     @       ������������������������       �        	             2@ K@lt �������������������������       �                     @    
   �       �                    '@�W�{�5�?�            �q@        �       �                     @��H�}�?             9@    ,   ������������������������       �                     @G   r   �       �                 ���A@      �?
             2@       �       �                    @ףp=
�?             $@    r   ������������������������       �                     �?    t   ������������������������       �                     "@   c   ������������������������       �                      @        �       �                 �?�@0Oex�I�?�            @p@    i   �       �                     @p� V�?=            �Y@    p   ������������������������       �                     @    )   �       �                    ?@@��8��?9             X@       �       �                   �8@@�z�G�?.             T@    l   �       �                    7@ ���J��?            �C@       ������������������������       �                     ?@   t   �       �                 `fF@      �?              @    a   �       �                 �&b@�q�q�?             @        ������������������������       �                      @   p   ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �D@   t   �       �                 �&B@      �?             0@   e   ������������������������       �        
             .@       ������������������������       �                     �?       �                          �?P��-�?h            �c@       �       �                     @0�I��8�?T             _@        �       �                    F@dP-���?!            �G@       �       �                   @D@������?            �B@   t   �       �                   �3@�#-���?            �A@       �       �                   �(@ȵHPS!�?             :@        �       �                   �5@$�q-�?             *@        �       �                    &@r�q��?             @        ������������������������       �                     �?    e   ������������������������       �                     @   n   ������������������������       �                     @    x   �       �                 �|�<@8�Z$���?
             *@    i   ������������������������       �                     @       �       �                   �A@�q�q�?             @   #   �       �                 �|�=@�q�q�?             @    .   ������������������������       �                     �?    t   �       �                    @@      �?              @    t   ������������������������       �                     �?       ������������������������       �                     �?       ������������������������       �                     @    a   ������������������������       �                     "@    r   ������������������������       �      �?              @       ������������������������       �                     $@       �                         @@@؇���X�?3            @S@       �       
                �|Y>@���*�?&             N@   _   �                       �!&B@�t����?!            �I@       �       �                   �1@�8��8��?             H@        ������������������������       �                     $@        �       �                   �2@�KM�]�?             C@        ������������������������       �                     �?    s   �       �                 ��) @�L���?            �B@    a   ������������������������       �                     4@   r   �                       @3�!@@�0�!��?             1@        �       �                 pf� @�q�q�?             @        ������������������������       �                     �?                               �|Y<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                �<@@4և���?             ,@       ������������������������       �                     &@                              �|Y=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @              	                   ;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                �?@X�<ݚ�?             "@        ������������������������       �                     @                              ��I @�q�q�?             @       ������������������������       ����Q��?             @        ������������������������       �                     �?        ������������������������       �                     1@        ������������������������       �                    �@@        �t�bh�h*h-K ��h/��R�(KMKK��h]�B       �{@     �p@      X@     @Y@     �Q@     �T@       @     �N@       @     �E@              6@       @      5@              @       @      0@       @                      0@              2@      Q@      6@      "@      (@       @      (@      @      @              @      @              @      @       @              �?      @              @      �?              �?             �M@      $@      2@             �D@      $@     �D@      "@      ;@      "@      .@      @      @       @              �?      @      �?      @              �?      �?      �?                      �?      &@       @      @       @       @               @       @      @              (@      @       @       @       @                       @      $@      @      @      @      @              @      @      @              ,@                      �?      :@      2@       @      .@       @      $@       @      �?              �?       @                      "@      @      @      �?      @              @      �?       @      �?                       @      @              2@      @      $@      @      $@      �?              �?      $@                       @       @             �u@     `d@      J@     �[@      *@      O@      &@      O@      @      H@              2@      @      >@      @      "@               @      @      @       @               @      @              @       @      �?       @                      �?              5@      @      ,@      @      ,@      @       @      @       @      �?      @              @      �?              @      @       @              �?      @              @      �?      �?      �?                      �?       @                      @      �?               @             �C@     �H@     �B@      =@      9@      6@              @      9@      1@      7@      .@      4@      .@      @              1@      .@      @      "@       @              �?      "@      �?      @              @      �?                      @      ,@      @      @              "@      @       @      @              @       @              @       @              �?      @      �?      @                      �?      @               @       @               @       @              (@      @              @      (@      �?       @              @      �?      @                      �?       @      4@      �?              �?      4@              $@      �?      $@      �?       @              �?      �?      �?      �?                      �?               @     �r@      J@     �G@      3@      *@      &@              @      *@      @      *@      @      &@      @       @              @      @              �?      @       @      @      �?       @              �?      �?      �?                      �?              �?       @       @      �?       @      �?      �?              �?      �?                       @      A@       @              @      A@      @      ?@      @      *@      @      "@              @      @       @               @      @       @      �?              �?       @                      @      2@              @             �o@     �@@      "@      0@              @      "@      "@      �?      "@      �?                      "@       @             `n@      1@     @Y@       @      @             �W@       @     �S@      �?      C@      �?      ?@              @      �?       @      �?       @                      �?      @             �D@              .@      �?      .@                      �?     �a@      .@     @[@      .@     �E@      @     �@@      @      @@      @      7@      @      (@      �?      @      �?              �?      @              @              &@       @      @              @       @      �?       @              �?      �?      �?      �?                      �?      @              "@              �?      �?      $@             �P@      &@     �H@      &@     �F@      @      F@      @      $@              A@      @              �?      A@      @      4@              ,@      @      �?       @              �?      �?      �?              �?      �?              *@      �?      &@               @      �?              �?       @              �?       @               @      �?              @      @              @      @       @      @       @      �?              1@             �@@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�ޡhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM%huh*h-K ��h/��R�(KM%��h|�B@I         �                 `f~I@�t����?�           8�@    @S@       S                    �?�����2�?�           h�@ 3��                          ��@V���#�?~            �g@     �Q@                        �|Y:@�IєX�?             1@     �?������������������������       �                     &@                                �&�@r�q��?             @        ������������������������       �                     �?      "@������������������������       �                     @      �?	                            @�.�8�?q            �e@        
                        ���*@�L#���?/            �P@                                `f�)@      �?             8@                                  �J@$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?                                  �B@"pc�
�?	             &@                                  :@�����H�?             "@                                   �?�q�q�?             @      @������������������������       �                     �?        ������������������������       �                      @     �[@������������������������       �                     @      2@                           D@      �?              @      @������������������������       �                     �?      �?������������������������       �                     �?      ,@                           E@ qP��B�?            �E@     @������������������������       �                     ?@                                    �?�8��8��?             (@        ������������������������       �                     @                                   �?r�q��?             @      6@������������������������       �                     �?      .@������������������������       �                     @               &                    @�k��V��?B            �Z@                %                    �?؇���X�?             ,@     @!       $                    @      �?              @      @"       #                 ��0@      �?             @       @������������������������       �                      @       @������������������������       �                      @      $@������������������������       �                     @      @������������������������       �                     @       @'       D                 03�1@�+Fi��?;             W@     @(       =                 �?�-@�ݜ����?'            �M@     :@)       ,                 �̌@�&!��?            �E@       @*       +                   �2@�z�G��?             $@      �?������������������������       �                     @      &@������������������������       �                     @       @-       .                   �1@:ɨ��?            �@@       @������������������������       �                     @      �?/       <                    �?PN��T'�?             ;@     @0       1                 `�X!@���y4F�?             3@       @������������������������       �                     @       @2       7                   �9@����X�?	             ,@     �?3       6                    4@      �?              @      @4       5                    �?�q�q�?             @      P@������������������������       �                      @      @������������������������       �                     �?       @������������������������       �                     @     �J@8       9                    �?      �?             @      $@������������������������       �                     �?      �?:       ;                    A@���Q��?             @       ������������������������       �                     @      0@������������������������       �                      @      @������������������������       �                      @      �?>       ?                   �0@      �?
             0@      @������������������������       �                     �?        @       C                   �;@��S�ۿ?	             .@       @A       B                    �?�q�q�?             @        ������������������������       �                     �?       @������������������������       �                      @      @������������������������       �                     (@        E       H                    @"pc�
�?            �@@       F       G                    �?�����?             5@        ������������������������       �                      @        ������������������������       �                     3@        I       J                 0C�7@�q�q�?             (@        ������������������������       �                     �?        K       L                    �?���!pc�?             &@        ������������������������       �                     @        M       N                    @      �?              @        ������������������������       �                      @        O       R                    @      �?             @       P       Q                   @C@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        T       m                 �?�@б΅t�?           �x@        U       l                    �?�wY;��?X             a@       V       k                 �Yu@     x�?S             `@       W       b                    �?���F6��?B            �X@        X       Y                 ���@�ݜ�?            �C@        ������������������������       �        	             .@        Z       [                   �6@�q�q�?             8@        ������������������������       �                      @        \       ]                  ��@��2(&�?             6@        ������������������������       �                     "@        ^       _                 �|Y=@�θ�?	             *@        ������������������������       �                     �?        `       a                 X��A@r�q��?             (@       ������������������������       �z�G�z�?             $@        ������������������������       �                      @        c       d                    7@(;L]n�?)             N@        ������������������������       �                     3@        e       j                 ��L@������?            �D@       f       g                 ���@�(\����?             D@        ������������������������       �                     5@        h       i                 ���@�}�+r��?             3@        ������������������������       �                     �?        ������������������������       �                     2@        ������������������������       �                     �?        ������������������������       �                     =@        ������������������������       �                      @        n       �                     �?|;�c� �?�            pp@        o       t                 �|�<@�q�q�?              H@        p       q                   �;@؇���X�?             @        ������������������������       �                      @        r       s                 `f�D@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        u       �                    �?���?            �D@       v       �                  �>@�d�����?             C@       w       �                    K@���Q��?             9@       x       �                   �G@���Q��?
             .@       y       ~                    �?���Q��?             $@        z       {                 `f&;@      �?             @        ������������������������       �                      @        |       }                 �|�=@      �?             @        ������������������������       �                     �?        ������������������������       �                     @               �                 03k:@      �?             @        �       �                   �D@      �?              @        ������������������������       �                     �? ��z�  ������������������������       �                     �? Wz�  ������������������������       �                      @��z�  ������������������������       �                     @ Xz�  �       �                 ���=@ףp=
�?             $@TMy� �������������������������       �                     "@�z�  ������������������������       �                     �?��z�  ������������������������       �        	             *@Sz�  ������������������������       �                     @ Uz�  �       �                    �?��ݼ��?�            �j@Qz�  �       �                     @�r����?W            �`@ Uz�  �       �                    �? "��u�?              I@ Vz�  ������������������������       �                     �?Uz�  �       �                    �?��<D�m�?            �H@Wz�  �       �                   �*@      �?             H@�z�  �       �                 `fF)@l��\��?             A@ �z�  ������������������������       �                     $@�z�  �       �                 �|�<@      �?             8@ ��z�  ������������������������       �                     *@�z�  �       �                   �F@���!pc�?             &@�z�  �       �                 �|�=@      �?             @ �z�  ������������������������       �                     �? �z�  �       �                    B@���Q��?             @ ��z�  ������������������������       �                      @ ��z�  ������������������������       ��q�q�?             @�z�  ������������������������       �                     @ �z�  ������������������������       �                     ,@�z�  ������������������������       �                     �?l�y�  �       �                    �?@�0�!��?7            @U@ Uz�  ������������������������       �                     @ Qz�  �       �                 @3�@����!�?4            �T@ Wz�  �       �                    :@�eP*L��?             &@ �z�  ������������������������       �                     @ �z�  �       �                   �?@����X�?             @ �z�  ������������������������       �                      @��z�  �       �                   �A@���Q��?             @ �z�  ������������������������       ��q�q�?             @��z�  ������������������������       �      �?              @�z�  �       �                    )@D��\��?-            �Q@ Tz�  ������������������������       �                     �?Vz�  �       �                 �|Y=@������?,            �Q@ ��z�  �       �                 ��Y @��a�n`�?             ?@ ��z�  �       �                   �3@      �?              @ �z�  ������������������������       �                     @ �z�  ������������������������       �                     @ Rz�  �       �                 `�X#@�㙢�c�?             7@Uz�  �       �                 ���"@���y4F�?             3@Wz�  �       �                 @�!@�r����?
             .@�z�  �       �                 pf� @�<ݚ�?             "@ ��z�  ������������������������       �                      @�z�  �       �                    8@����X�?             @Tz�  ������������������������       �                     @ Vz�  ������������������������       �                      @ ��z�  ������������������������       �                     @ Uz�  �       �                   �<@      �?             @Wz�  ������������������������       �                      @j�y�  ������������������������       �                      @ ��z�  ������������������������       �                     @��z�  �       �                   �?@�7��?            �C@�z�  �       �                 ��) @���}<S�?             7@Vz�  ������������������������       �                     ,@ Wz�  �       �                 �|�=@�<ݚ�?             "@�z�  �       �                 pf� @      �?              @ Qz�  ������������������������       �                     �?Wz�  ������������������������       �                     @�z�  ������������������������       �                     �? �z�  ������������������������       �        	             0@�z�  �       �                    �?�z�G��?5             T@ �z�  �       �                 �2@�n_Y�K�?             *@�z�  �       �                 �|�;@�����H�?             "@Uz�  �       �                 �&�)@      �?             @ l�y�  ������������������������       �                      @Wz�  �       �                    �?      �?              @ Wz�  ������������������������       �                     �?Sz�  ������������������������       �                     �? �z�  ������������������������       �                     @�z�  ������������������������       �                     @Wz�  �       �                    �?���}D�?-            �P@ �z�  �       �                    �? ��WV�?             :@ �z�  ������������������������       �                     @ �z�  �       �                    6@�nkK�?             7@ �z�  ������������������������       �                     �? Tz�  ������������������������       �                     6@ Vz�  �       �                    @��]�T��?            �D@��z�  �       �                    �?\�Uo��?             C@ �z�  ������������������������       �                      @��z�  �       �                    @�q�q�?             B@�z�  �       �                 03{3@�q�����?             9@ �z�  �       �                     @z�G�z�?             $@ ��z�  �       �                    *@z�G�z�?             @ Wz�  ������������������������       �                     �?�z�  ������������������������       �                     @��z�  �       �                   �5@z�G�z�?             @Uz�  ������������������������       �                     @ Wz�  ������������������������       �                     �? �z�  �       �                 �̌4@�q�q�?             .@ �z�  ������������������������       �                     @ �z�  �       �                    �?�q�q�?             (@m�y�  �       �                    :@�z�G��?             $@�z�  �       �                     @      �?             @ �z�  ������������������������       �                      @�z�  �       �                    +@      �?              @ �z�  ������������������������       �                     �? i�y�  ������������������������       �                     �?    s   ������������������������       �                     @   #   ������������������������       �                      @    k   �       �                    �?"pc�
�?             &@    g   ������������������������       �                     @   i   �       �                 pf�C@�q�q�?             @    b   �       �                    @�q�q�?             @        ������������������������       �                      @   p   ������������������������       �                     �?   t   ������������������������       �                     @   f   ������������������������       �                     @    g   �       �                    �?ƆQ����?P            �^@   _   �       �                  "�b@pY���D�?0            �S@   l   ������������������������       �        %            �M@        �       �                    �?ףp=
�?             4@   s   ������������������������       �                     $@    a   �       �                    $@z�G�z�?             $@        ������������������������       �                      @   a   ������������������������       �                      @        �                           @�&!��?             �E@       �                          �?p�ݯ��?             C@   a   �                           �?b�2�tk�?             B@   f   �       	                �UwR@���Q��?            �A@    e   �                          �?�<ݚ�?             2@                                  �?���Q��?             @    t   ������������������������       �                      @                              ��UO@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                                �C@$�q-�?             *@        ������������������������       �                     @                                 F@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        
                         �?j���� �?             1@                                 �?      �?              @                                �?؇���X�?             @                                �9@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?                                 �?X�<ݚ�?             "@                                �?z�G�z�?             @                              �̾w@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                 �?      �?             @                                =@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @              $                p�O@���Q��?             @              #                   >@      �?             @       !      "                   ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �t�b�[     h�h*h-K ��h/��R�(KM%KK��h]�BP       �z@     �q@     �x@      h@      O@      `@      �?      0@              &@      �?      @      �?                      @     �N@      \@      @     �O@      @      5@      �?      (@              (@      �?               @      "@      �?       @      �?       @      �?                       @              @      �?      �?      �?                      �?      �?      E@              ?@      �?      &@              @      �?      @      �?                      @     �L@     �H@       @      (@       @      @       @       @               @       @                      @              @     �K@     �B@      <@      ?@      :@      1@      @      @      @                      @      7@      $@              @      7@      @      .@      @      @              $@      @      @      �?       @      �?       @                      �?      @              @      @      �?               @      @              @       @               @               @      ,@      �?              �?      ,@      �?       @      �?                       @              (@      ;@      @      3@       @               @      3@               @      @              �?       @      @      @              @      @       @              @      @       @      @              @       @              �?             �t@     @P@      `@      @     @^@      @      W@      @      A@      @      .@              3@      @               @      3@      @      "@              $@      @              �?      $@       @       @       @       @              M@       @      3@             �C@       @     �C@      �?      5@              2@      �?              �?      2@                      �?      =@               @             �i@      M@      @@      0@      �?      @               @      �?      @              @      �?              ?@      $@      <@      $@      .@      $@      @      "@      @      @      @      @               @      @      �?              �?      @              @      �?      �?      �?              �?      �?               @                      @      "@      �?      "@                      �?      *@              @             �e@      E@     @]@      2@     �G@      @      �?              G@      @     �F@      @      ?@      @      $@              5@      @      *@               @      @      @      @              �?      @       @       @              �?       @      @              ,@              �?             �Q@      .@      @             �P@      .@      @      @      @               @      @               @       @      @      �?       @      �?      �?     �N@      $@              �?     �N@      "@      8@      @      @      @              @      @              3@      @      .@      @      *@       @      @       @       @              @       @      @                       @      @               @       @       @                       @      @             �B@       @      5@       @      ,@              @       @      @      �?              �?      @                      �?      0@              L@      8@      @       @      �?       @      �?      @               @      �?      �?      �?                      �?              @      @             �I@      0@      9@      �?      @              6@      �?              �?      6@              :@      .@      7@      .@       @              5@      .@      (@      *@       @       @      �?      @      �?                      @      �?      @              @      �?              $@      @      @              @      @      @      @      �?      @               @      �?      �?              �?      �?              @                       @      "@       @      @              @       @      �?       @               @      �?              @              @              <@     �W@       @     @S@             �M@       @      2@              $@       @       @       @                       @      :@      1@      8@      ,@      6@      ,@      5@      ,@      ,@      @       @      @               @       @      �?       @                      �?      (@      �?      @              @      �?              �?      @              @      $@       @      @      �?      @      �?       @      �?                       @              @      �?              @      @      @      �?      �?      �?      �?                      �?      @              �?      @      �?      �?              �?      �?                       @      �?               @               @      @      �?      @      �?      �?              �?      �?                       @      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJQY%hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtK�huh*h-K ��h/��R�(KK���h|�B�?                             @��ϙLq�?�           8�@               	                    @     ��?             @@                                  @��.k���?             1@���                             �?ףp=
�?             $@      @                             @      �?              @      @������������������������       �                     �?      E@������������������������       �                     �?      @������������������������       �                      @      (@������������������������       �                     @      �?
                           �?��S�ۿ?
             .@     @������������������������       �                     $@       @                           @z�G�z�?             @       @������������������������       �                     @                                   �?      �?              @       @������������������������       �                     �?        ������������������������       �                     �?      @       �                 `fK@�ĸۦ��?�           8�@     @       Q                    �?��J��?r           @�@      @       "                     @Z�2�t��?h            �d@      @       !                    �?0)RH'�?(            @Q@      @                          �*@�q�q��?             H@       @                           B@���Q��?             4@     @                          �9@      �?	             0@      @                          �'@z�G�z�?             @       @������������������������       �                     �?       @������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     @     @U@                        ���;@ �Cc}�?             <@       ������������������������       �                     6@     �I@                         X��C@      �?             @     &@������������������������       �                     @        ������������������������       �                     @ ���  ������������������������       �                     5@�8��  #       0                 pF @�W*��?@            @X@ ���  $       /                    �?��hJ,�?             A@���  %       .                 X��B@<���D�?            �@@���  &       '                   �6@     ��?             @@ >��  ������������������������       �                     .@ ��  (       )                   �8@@�0�!��?             1@ ��  ������������������������       �                      @0��  *       -                 ���@��S�ۿ?             .@ ��  +       ,                 �Y�@      �?             @ ��  ������������������������       �                     @ ���  ������������������������       �                     �?     �?������������������������       �        	             &@���  ������������������������       �                     �?��  ������������������������       �                     �? ���  1       N                 03�7@����X�?+            �O@N��  2       K                    �?�D����?             E@���  3       F                    �?p�ݯ��?             C@     @4       ?                 ��.@     ��?             @@���  5       >                    �?�J�4�?             9@���  6       ;                 �&�%@������?             1@���  7       :                 `��!@ףp=
�?             $@ ���  8       9                 `�X!@      �?             @��  ������������������������       �                     @ ���  ������������������������       �                     �? ���  ������������������������       �                     @0��  <       =                 ���*@և���X�?             @ <��  ������������������������       �                     @���  ������������������������       �                     @ ���  ������������������������       �                      @b��  @       A                    �?؇���X�?             @ ��  ������������������������       �                     @      �?B       C                 03�1@      �?             @      �?������������������������       �                      @      @D       E                    �?      �?              @      @������������������������       �                     �?      �?������������������������       �                     �?      @G       J                    @�q�q�?             @      @H       I                   �4@���Q��?             @      @������������������������       �                      @       @������������������������       �                     @        ������������������������       �                     �?        L       M                 �|Y=@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        O       P                    �?���N8�?             5@        ������������������������       �                     �?        ������������������������       �                     4@        R       �                   �J@T�1!�}�?
            z@       S       \                   �2@      �?�            �x@        T       [                 �&@������?             B@        U       V                    �?�X�<ݺ?             2@       ������������������������       �                     $@        W       Z                    �?      �?              @        X       Y                  �K"@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     2@        ]       x                     �?4�<����?�            @v@        ^       e                 �|�<@��J�fj�?            �B@        _       `                    7@      �?              @        ������������������������       �                     �?        a       b                 `f�D@؇���X�?             @       ������������������������       �                     @        c       d                 ��I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        f       w                   �G@J�8���?             =@       g       r                 �TA@@l��
I��?             ;@       h       m                 ���=@j���� �?             1@       i       l                 ��";@"pc�
�?
             &@       j       k                 ��:@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        n       o                  �>@r�q��?             @        ������������������������       �                     @        p       q                  �>@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        s       t                   �C@ףp=
�?             $@       ������������������������       �                     @        u       v                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        y       �                    �?0�\>��?�            �s@       z       �                   @E@�u����?�             q@       {       �                    �?Ǖi�7�?�            0p@       |       �                     @X�EQ]N�?�             p@        }       ~                    �?���c���?             J@        ������������������������       �                     @               �                   @D@؇���X�?            �H@       �       �                 `fF)@�����H�?            �F@        �       �                    5@���7�?             6@ ��z�  ������������������������       �                     �? Wz�  ������������������������       �                     5@��z�  �       �                 �|�<@�㙢�c�?             7@ Xz�  ������������������������       �                      @TMy� ��       �                   �3@������?             .@�z�  �       �                   �A@�	j*D�?             *@�z�  �       �                    @@      �?              @Sz�  �       �                 �|�=@      �?             @ Uz�  ������������������������       �                     �?Qz�  ������������������������       �                     @ Uz�  ������������������������       �      �?             @ Vz�  ������������������������       �                     @Uz�  ������������������������       �                      @Wz�  ������������������������       �      �?             @�z�  �       �                 �Y�@�"�_*d�?�            �i@ �z�  �       �                   �8@���y4F�?             C@ �z�  �       �                   �3@���|���?             &@ ��z�  ������������������������       �                     @�z�  �       �                    5@      �?              @ �z�  �       �                    �?�q�q�?             @ �z�  ������������������������       �                      @ �z�  ������������������������       �                     �? ��z�  ������������������������       �                     @ ��z�  �       �                 ���@ 7���B�?             ;@�z�  ������������������������       �                     6@ �z�  ������������������������       �z�G�z�?             @�z�  �       �                 �?�@4և����?k             e@l�y�  �       �                 �?$@x��B�R�?9            �V@ Uz�  �       �                    ;@�8��8��?             B@ Qz�  ������������������������       �                     *@ Wz�  �       �                  s�@�LQ�1	�?             7@ �z�  ������������������������       �                     @ �z�  �       �                    �?     ��?             0@�z�  �       �                 �|Y=@"pc�
�?	             &@ ��z�  ������������������������       �                     �? �z�  �       �                 X��A@ףp=
�?             $@��z�  ������������������������       ������H�?             "@�z�  ������������������������       �                     �? Tz�  �       �                 �|Y>@z�G�z�?             @ Vz�  ������������������������       �      �?              @ ��z�  ������������������������       �                     @ ��z�  ������������������������       �                    �K@ �z�  �       �                    �?� ���?2            @S@ �z�  ������������������������       �                     @ Rz�  �       �                   @C@�MI8d�?/            �R@Uz�  �       �                   �3@؇���X�?,            �Q@ Wz�  ������������������������       ����Q��?             @�z�  �       �                 ��) @�?�<��?*            @P@��z�  �       �                   �>@��(\���?             D@�z�  ������������������������       �                     =@Tz�  �       �                   �@@���!pc�?             &@Vz�  �       �                   �?@      �?             @ ��z�  ������������������������       �                     �? Uz�  ������������������������       ����Q��?             @Wz�  ������������������������       �                     @j�y�  �       �                 �|�>@z�G�z�?             9@��z�  �       �                   �8@      �?             4@ ��z�  ������������������������       �                     @�z�  �       �                 0S%"@     ��?             0@ Vz�  �       �                 �|Y<@���Q��?             @ Wz�  ������������������������       �                      @�z�  �       �                 pf� @�q�q�?             @ Qz�  ������������������������       �                     �?Wz�  ������������������������       �                      @�z�  �       �                   �<@"pc�
�?             &@ �z�  ������������������������       �                     @�z�  �       �                 �|Y=@���Q��?             @ �z�  �       �                 ���"@�q�q�?             @ �z�  ������������������������       �                     �?Uz�  ������������������������       �                      @ l�y�  ������������������������       �                      @Wz�  ������������������������       �                     @ Wz�  �       �                   @D@      �?             @Sz�  �       �                 ��	0@�q�q�?             @ �z�  ������������������������       �                      @�z�  ������������������������       �                     �?Wz�  ������������������������       �                     �? �z�  ������������������������       �                     �? �z�  ������������������������       �                     .@ �z�  �       �                 ��.@`Ӹ����?            �F@ �z�  �       �                    �?r�q��?	             (@Tz�  �       �                     @�C��2(�?             &@ Vz�  ������������������������       �                     �?��z�  �       �                    5@ףp=
�?             $@ �z�  ������������������������       �                     �?��z�  ������������������������       �                     "@�z�  ������������������������       �                     �? �z�  ������������������������       �                    �@@ ��z�  ������������������������       �                     :@ Wz�  �       �                    �?�"�q��?A            �W@�z�  �       �                    �?�}�+r��?'            �L@��z�  ������������������������       �                     =@Uz�  �       �                    @ �Cc}�?             <@Wz�  ������������������������       �                     9@ �z�  ������������������������       �                     @ �z�  �       �                    �?p�ݯ��?             C@�z�  �       �                 X�,@@��Q��?             4@m�y�  �       �                  �}S@      �?             $@ �z�  ������������������������       �                     @ �z�  �       �                    �?r�q��?             @�z�  ������������������������       �                     @ �z�  �       �                   �5@      �?              @ i�y�  ������������������������       �                     �?    s   ������������������������       �                     �?   #   �       �                    �?z�G�z�?             $@   k   �       �                   @H@�����H�?             "@   g   ������������������������       �                     @   i   �       �                   �T@�q�q�?             @    b   ������������������������       �                      @        ������������������������       �                     �?   p   ������������������������       �                     �?   t   �       �                     @b�2�tk�?             2@   f   �       �                     �?      �?	             (@   g   �       �                 �|Y>@�eP*L��?             &@    _   ������������������������       �                     �?   l   �       �                    �?���Q��?             $@       �       �                 03�U@      �?              @   s   �       �                    C@�q�q�?             @    a   ������������������������       �                     �?        ������������������������       �                      @   a   ������������������������       �                     @        ������������������������       �                      @       ������������������������       �                     �?   a   �       �                    @r�q��?             @   f   ������������������������       �                     @    e   ������������������������       �                     �?        �t�bh�h*h-K ��h/��R�(KK�KK��h]�B�       �|@     �o@      "@      7@       @      "@      �?      "@      �?      �?      �?                      �?               @      @              �?      ,@              $@      �?      @              @      �?      �?      �?                      �?     �{@      m@     �z@     @c@     �N@     @Z@      &@      M@      &@     �B@       @      (@      @      (@      @      �?              �?      @                      &@      @              @      9@              6@      @      @              @      @                      5@      I@     �G@      @      =@      @      =@      @      =@              .@      @      ,@       @              �?      ,@      �?      @              @      �?                      &@      �?              �?             �F@      2@      9@      1@      8@      ,@      6@      $@      5@      @      *@      @      "@      �?      @      �?      @                      �?      @              @      @              @      @               @              �?      @              @      �?      @               @      �?      �?      �?                      �?       @      @       @      @       @                      @              �?      �?      @              @      �?              4@      �?              �?      4@             w@     �H@     pu@     �H@     �A@      �?      1@      �?      $@              @      �?      @      �?      @                      �?      @              2@             @s@      H@      5@      0@       @      @      �?              �?      @              @      �?      �?      �?                      �?      3@      $@      3@       @      $@      @      "@       @      @       @      @                       @      @              �?      @              @      �?       @      �?                       @      "@      �?      @              @      �?      @                      �?               @     �q@      @@     �n@      >@     �l@      >@     �l@      >@     �F@      @      @              E@      @      D@      @      5@      �?              �?      5@              3@      @       @              &@      @      "@      @      @      @      @      �?              �?      @              �?      @      @               @               @       @     �f@      7@      >@       @      @      @      @              �?      @      �?       @               @      �?                      @      :@      �?      6@              @      �?      c@      .@      V@      @     �@@      @      *@              4@      @      @              *@      @      "@       @              �?      "@      �?       @      �?      �?              @      �?      �?      �?      @             �K@             @P@      (@      @              O@      (@      N@      $@      @       @     �L@       @     �B@      @      =@               @      @      @      @              �?      @       @      @              4@      @      .@      @      @              &@      @       @      @               @       @      �?              �?       @              "@       @      @              @       @      �?       @      �?                       @       @              @               @       @      �?       @               @      �?              �?              �?              .@             �E@       @      $@       @      $@      �?      �?              "@      �?              �?      "@                      �?     �@@              :@              1@     �S@      @      K@              =@      @      9@              9@      @              ,@      8@      @      *@      @      @              @      @      �?      @              �?      �?      �?                      �?       @       @      �?       @              @      �?       @               @      �?              �?              @      &@      @      @      @      @      �?              @      @       @      @       @      �?              �?       @                      @       @              �?              �?      @              @      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ��fbhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM5huh*h-K ��h/��R�(KM5��h|�B@M         F                    �?�u����?�           8�@                                   �?sYi9��?O            `a@                                    @\#r��?"            �N@���                            �H@��<b�ƥ?             G@     @������������������������       �                     E@      M@                           J@      �?             @      �?������������������������       �                     �?        ������������������������       �                     @      @	                           �?�q�q�?
             .@       
                           �?X�Cc�?	             ,@                                �&�)@և���X�?             @      4@������������������������       �                     @      @������������������������       �                     @      ,@                        `�@1@����X�?             @                                  @      �?             @      �?������������������������       �                      @     �?������������������������       �                      @      �?������������������������       �                     @      @������������������������       �                     �?      @       E                 �U�X@�θ�?-            �S@     �?       D                  �	U@��R[s�?*            �Q@     �?       C                    �?��ga�=�?(            �P@     �?       <                 ��<J@�'�`d�?'            �P@              9                    �?&y�X���?#             M@              6                    �?r�����?             �J@              5                 p�i@@��k=.��?            �G@     @       2                   `A@�I�w�"�?             C@      @       1                 �|�=@"pc�
�?            �@@      @                             �?d}h���?             <@                                0C�<@      �?              @       @������������������������       �                     �?      >@������������������������       �                     �?      @!       (                    ;@���B���?             :@      @"       '                 ���@�8��8��?             (@      @#       $                 ��y@؇���X�?             @       @������������������������       �                     �?      $@%       &                   �7@r�q��?             @      @������������������������       �                     �?       @������������������������       �                     @     @������������������������       �                     @     :@)       *                 �|Y=@����X�?	             ,@       @������������������������       �                     �?      �?+       ,                     @�θ�?             *@      &@������������������������       �                     �?       @-       0                   @@      �?             (@      @.       /                 ���@      �?              @      �?������������������������       �                     �?     @������������������������       �և���X�?             @       @������������������������       �                     @       @������������������������       �                     @     �?3       4                      @���Q��?             @      @������������������������       �                     @      P@������������������������       �                      @      @������������������������       �                     "@       @7       8                 �&�)@r�q��?             @     �J@������������������������       �                     �?      $@������������������������       �                     @      �?:       ;                ��k/@z�G�z�?             @        ������������������������       �                     �?      0@������������������������       �                     @      @=       B                 ���Q@      �?              @     �?>       A                    �?      �?             @     @?       @                    F@      �?              @        ������������������������       �                     �?       @������������������������       �                     �?        ������������������������       �                      @       @������������������������       �                     @      @������������������������       �                     �?        ������������������������       �                     @       ������������������������       �                      @        G                          �?��s�ɝ�?t           ��@       H       �                    �?>4և���?"            |@       I       z                    �?������?�            �w@        J       g                   �9@z�G�z�?2            �R@        K       `                   �6@�û��|�?             7@       L       _                 8#B2@������?             1@       M       N                   �1@���|���?
             &@        ������������������������       �                     �?        O       X                   �4@���Q��?	             $@       P       Q                    �?      �?             @        ������������������������       �                     �?        R       W                    3@���Q��?             @       S       T                 P��@      �?             @        ������������������������       �                     �?        U       V                 ��!@�q�q�?             @        ������������������������       �                      @       ������������������������       �                     �?        ������������������������       �                     �?        Y       Z                     @      �?             @        ������������������������       �                     �?        [       \                    �?�q�q�?             @        ������������������������       �                     �?        ]       ^                 pF�!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @       a       b                     @r�q��?             @        ������������������������       �                     �?        c       f                    8@z�G�z�?             @       d       e                 @3�@�q�q�?             @        ������������������������       �                     �?       ������������������������       �                      @        ������������������������       �                      @        h       i                    �?ȵHPS!�?!             J@        ������������������������       �                     $@        j       w                     @؇���X�?             E@       k       n                 `f&'@ >�֕�?            �A@        l       m                   �E@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        o       p                     �?�g�y��?             ?@        ������������������������       �                     *@        q       r                   �B@�X�<ݺ?             2@       ������������������������       �                     "@       s       v                   �*@�����H�?             "@        t       u                    D@      �?             @        ������������������������       �                     �?       ������������������������       �                     @       ������������������������       �                     @       x       y                 �|�;@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        {       �                 ��$:@�Qb��?�            �r@       |       �                   @@@������?�            0p@       }       �                   �>@$�3c�s�?v            �g@       ~       �                 @3�@��I�� �?o            `f@              �                 �|Y=@��<D�m�?;            �X@        �       �                 ��@      �?             D@       �       �                  ��@z�G�z�?             9@��z�  �       �                    �?�C��2(�?             6@ Wz�  ������������������������       �                     �?��z�  �       �                    7@�����?             5@Xz�  ������������������������       �                     (@TMy� ��       �                 ���@�<ݚ�?             "@ �z�  �       �                 �&b@�q�q�?             @ �z�  ������������������������       �                     �?Sz�  ������������������������       �                      @ Uz�  ������������������������       �                     @Qz�  ������������������������       �                     @ Uz�  ������������������������       �                     .@ Vz�  �       �                 �|�=@ _�@�Y�?             M@Uz�  �       �                     @@3����?             K@ Wz�  ������������������������       �                     &@�z�  �       �                 ��@ qP��B�?            �E@�z�  ������������������������       �                     6@ �z�  �       �                 �Y5@���N8�?
             5@ ��z�  ������������������������       �z�G�z�?             @�z�  ������������������������       �                     0@ �z�  ������������������������       �                     @ �z�  �       �                   �3@�
��P�?4            @T@ �z�  �       �                   �2@�d�����?             3@��z�  �       �                 ��Y @ףp=
�?             $@ ��z�  �       �                    1@      �?              @ �z�  ������������������������       �                     �? �z�  ������������������������       �                     �?�z�  ������������������������       �                      @l�y�  �       �                 ���$@X�<ݚ�?             "@Uz�  �       �                 0S5 @����X�?             @ Qz�  ������������������������       ��q�q�?             @ Wz�  ������������������������       �                     @ �z�  ������������������������       �                      @ �z�  �       �                    �?��a�n`�?(             O@ �z�  ������������������������       �                     �? ��z�  �       �                 ��) @\#r��?'            �N@ �z�  ������������������������       �                     6@��z�  �       �                    :@8�Z$���?            �C@ �z�  ������������������������       �                     .@ Tz�  �       �                     @      �?             8@ Vz�  �       �                 �|Y<@�8��8��?             (@ ��z�  ������������������������       �                     @ ��z�  �       �                     �?؇���X�?             @ �z�  ������������������������       �                      @ �z�  �       �                 �|�=@z�G�z�?             @ Rz�  ������������������������       �                     �?Uz�  ������������������������       �                     @ Wz�  �       �                 0S%"@�q�q�?             (@ �z�  �       �                 pf� @z�G�z�?             @ ��z�  ������������������������       �                      @�z�  �       �                 �|Y<@�q�q�?             @ Tz�  ������������������������       �                      @Vz�  ������������������������       �                     �? ��z�  �       �                 �|�=@؇���X�?             @Uz�  ������������������������       �                     @Wz�  ������������������������       �                     �?j�y�  �       �                 �&B@X�<ݚ�?             "@ ��z�  ������������������������       �                     �? ��z�  �       �                   �@      �?              @ �z�  ������������������������       �                     @ Vz�  �       �                 �?�@���Q��?             @ Wz�  ������������������������       �                     �?�z�  �       �                 ��I @      �?             @Qz�  �       �                   �?@�q�q�?             @ Wz�  ������������������������       �                     �?�z�  ������������������������       �      �?              @ �z�  ������������������������       �                     �?�z�  �       �                   @E@�J�T�?-            �Q@�z�  �       �                 �?�@�X�<ݺ?             B@ �z�  ������������������������       �        
             1@Uz�  �       �                 @3�@�KM�]�?             3@ l�y�  ������������������������       ��q�q�?             @Wz�  �       �                   @D@      �?             0@Wz�  ������������������������       �                     ,@Sz�  �       �                     @      �?              @ �z�  ������������������������       �                     �?�z�  ������������������������       �                     �?Wz�  ������������������������       �                    �A@ �z�  �       �                     �?X��ʑ��?            �E@�z�  �       �                 ��yC@j���� �?             A@�z�  �       �                   �A@����X�?             <@�z�  �       �                 �T!@@�q�q�?             8@Tz�  �       �                   �J@���!pc�?             6@Vz�  �       �                 `fF<@�t����?	             1@��z�  �       �                 �|�?@$�q-�?             *@ �z�  ������������������������       �                     �?��z�  ������������������������       �                     (@�z�  �       �                   @>@      �?             @ �z�  ������������������������       �                     �? ��z�  ������������������������       �                     @ Wz�  �       �                 `fF<@z�G�z�?             @�z�  ������������������������       �                     @��z�  ������������������������       �                     �?Uz�  ������������������������       �                      @Wz�  ������������������������       �                     @ �z�  ������������������������       �                     @ �z�  �       �                    ;@�<ݚ�?             "@ �z�  �       �                 ��?P@�q�q�?             @ m�y�  ������������������������       �                      @ �z�  ������������������������       �                     �? �z�  ������������������������       �                     @�z�  �       �                   �:@DX�\��?3            �Q@ �z�  �       �                    �?��2(&�?             6@i�y�  �       �                     @     ��?             0@    s   �       �                    2@����X�?             @    #   ������������������������       �                     �?   k   �       �                     �?r�q��?             @    g   ������������������������       �                      @   i   �       �                    �?      �?             @    b   ������������������������       �                     �?        ������������������������       �                     @   p   �       �                   �!@�����H�?             "@    t   �       �                 ��Y@      �?             @    f   ������������������������       �                     @   g   ������������������������       �                     �?    _   ������������������������       �                     @   l   ������������������������       �                     @       �       �                    �?Rg��J��?%            �H@    s   �       �                   @C@���|���?             &@   a   �       �                    �?�z�G��?             $@       ������������������������       �                     @   a   ������������������������       �                     @        ������������������������       �                     �?       �                           @      �?             C@   a   �                         @D@��}*_��?             ;@   f   �                           �?�<ݚ�?             2@   e   �                       �|Y=@r�q��?	             (@                               ���M@      �?              @    t   ������������������������       �                     �?        ������������������������       �                     �?                                 �?ףp=
�?             $@       ������������������������       �                     @                              `f�K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                �@@�q�q�?             @       	      
                  �<@z�G�z�?             @        ������������������������       �                     �?                                �7@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                                  �?�q�q�?             "@                             �CdQ@      �?              @        ������������������������       �                     @                                 �?���Q��?             @        ������������������������       �                      @                              ��#[@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?                                 �?"pc�
�?             &@                              ���.@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @              (                    @�^�����?R             _@                                 �? i���t�?$            �H@       ������������������������       �                     C@               !                   �?�eP*L��?             &@        ������������������������       �                     �?        "      '                   �?���Q��?             $@       #      $                    �?X�<ݚ�?             "@        ������������������������       �                      @        %      &                   :@����X�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        )      4                   �?��n�?.            �R@        *      +                  �7@���Q��?            �A@        ������������������������       �                     (@        ,      1                ��T?@���}<S�?             7@       -      0                   @@�}�+r��?             3@        .      /                �|Y>@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             ,@        2      3                ���A@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     D@        �t�bh�h*h-K ��h/��R�(KM5KK��h]�BP       �{@     �p@     �P@     @R@      @     �K@      �?     �F@              E@      �?      @      �?                      @      @      $@      @      "@      @      @              @      @               @      @       @       @               @       @                      @              �?      N@      2@      J@      2@      J@      .@      J@      ,@     �G@      &@     �E@      $@      C@      "@      =@      "@      ;@      @      6@      @      �?      �?      �?                      �?      5@      @      &@      �?      @      �?      �?              @      �?              �?      @              @              $@      @              �?      $@      @      �?              "@      @      @      @      �?              @      @      @              @               @      @              @       @              "@              @      �?              �?      @              @      �?              �?      @              @      @      �?      @      �?      �?              �?      �?                       @      @                      �?              @       @             �w@      h@     �s@     �`@     �p@     �Z@      .@      N@      "@      ,@      @      *@      @      @              �?      @      @      @      @              �?      @       @       @       @              �?       @      �?       @                      �?      �?              �?      @              �?      �?       @              �?      �?      �?              �?      �?                      @      @      �?      �?              @      �?       @      �?              �?       @               @              @      G@              $@      @      B@       @     �@@      �?      @              @      �?              �?      >@              *@      �?      1@              "@      �?       @      �?      @      �?                      @              @      @      @              @      @              p@      G@     `m@      8@     �d@      6@     @d@      1@      W@      @     �A@      @      4@      @      4@       @      �?              3@       @      (@              @       @      �?       @      �?                       @      @                      @      .@             �L@      �?     �J@      �?      &@              E@      �?      6@              4@      �?      @      �?      0@              @             �Q@      &@      ,@      @      "@      �?      �?      �?      �?                      �?       @              @      @      @       @      �?       @      @                       @      L@      @      �?             �K@      @      6@             �@@      @      .@              2@      @      &@      �?      @              @      �?       @              @      �?              �?      @              @      @      �?      @               @      �?       @               @      �?              @      �?      @                      �?      @      @      �?              @      @              @      @       @      �?               @       @      �?       @              �?      �?      �?      �?             @Q@       @      A@       @      1@              1@       @       @      �?      .@      �?      ,@              �?      �?              �?      �?             �A@              5@      6@      ,@      4@       @      4@       @      0@      @      0@       @      .@      �?      (@      �?                      (@      �?      @      �?                      @      @      �?      @                      �?       @                      @      @              @       @      �?       @               @      �?              @              E@      =@      3@      @      *@      @      @       @              �?      @      �?       @              @      �?              �?      @               @      �?      @      �?      @                      �?      @              @              7@      :@      @      @      @      @              @      @              �?              3@      3@      $@      1@      @      ,@       @      $@      �?      �?              �?      �?              �?      "@              @      �?       @      �?                       @       @      @      �?      @              �?      �?      @      �?                      @      �?              @      @      @      @      @               @      @               @       @      �?       @                      �?      �?              "@       @      �?       @      �?                       @       @             �P@      M@      @      F@              C@      @      @      �?              @      @      @      @       @               @      @              @       @                      �?     �N@      ,@      5@      ,@              (@      5@       @      2@      �?      @      �?      @                      �?      ,@              @      �?              �?      @              D@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ$�phG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtK�huh*h-K ��h/��R�(KK���h|�B@?         .                   �3@�L*�<�?�           8�@               +                    @b�L�4��?P            �`@                                  �?�Sb(�	�?A             [@     �Q@                           �?���.�6�?             G@      �?������������������������       �        
             2@      2@                            @ �Cc}�?             <@     &@������������������������       �                     2@      @       	                    @�z�G��?             $@      �?������������������������       �                     @        
                           �?      �?             @                                  �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @                                �?�@�g�y��?#             O@        ������������������������       �                     ,@                                   �?      �?             H@      �?������������������������       �                      @      @                            �?�LQ�1	�?             G@      @                           �?և���X�?             <@     �?                            @      �?
             8@      �?                          �2@      �?             @      �?������������������������       �                      @                                 �'@      �?             @        ������������������������       �                     @       ������������������������       �                     �?     @                        ��Y @      �?             2@      @                           1@ףp=
�?             $@       @������������������������       �      �?             @        ������������������������       �                     @       @������������������������       �                      @      >@������������������������       �                     @      @!       "                    �?�<ݚ�?             2@      @������������������������       �                      @      @#       $                 03{3@      �?             0@        ������������������������       �                     $@      @%       *                    �?�q�q�?             @       &       )                    �?���Q��?             @       '       (                    7@      �?             @      @������������������������       �                      @        ������������������������       �                      @      @������������������������       �                     �?       @������������������������       �                     �?        ,       -                   -@$�q-�?             :@       @������������������������       �                      @      @������������������������       �                     8@    �A@/       p                    �?B�����?_           �@      :@0       A                     @tHN�?q             f@      @1       >                   @L@X'"7��?H             [@       2       3                    �?T��,��?D            @Y@      "@������������������������       �                     A@       @4       =                    �?�����?-            �P@       5       6                   �B@@4և���?             E@     @������������������������       �                     =@      &@7       8                   @C@�θ�?	             *@       @������������������������       �                     �?        9       :                     �?r�q��?             (@       @������������������������       �                     @       ;       <                    �?����X�?             @     @������������������������       �                     @     @������������������������       �                      @      �?������������������������       �                     9@       ?       @                   �L@����X�?             @      @������������������������       �                      @     @������������������������       �                     @        B       m                    @\X��t�?)            @Q@      @C       l                 03�:@p�EG/��?%            �O@     @D       S                    �?d��0u��?"             N@        E       R                    �?������?             >@       F       Q                 ��.@l��
I��?             ;@       G       H                 �|Y=@X�<ݚ�?	             2@        ������������������������       �                     �?       I       N                    �?��.k���?             1@        J       M                    �?�<ݚ�?             "@       K       L                 X�x&@�q�q�?             @        ������������������������       �                      @       ������������������������       �                     @        ������������������������       �                     @        O       P                 �&�@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@       ������������������������       �                     @        T       k                   @B@��S���?             >@       U       f                    �?�5��?             ;@       V       ]                    �?      �?             4@       W       Z                 ��� @��
ц��?             *@       X       Y                   �9@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        [       \                    ;@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ^       _                 ���)@և���X�?             @        ������������������������       �                      @        `       e                 03�1@���Q��?             @       a       d                   �0@      �?             @       b       c                 �|�;@      �?              @        ������������������������       �                     �?       ������������������������       �                     �?        ������������������������       �                      @       ������������������������       �                     �?        g       h                    �?؇���X�?             @        ������������������������       �                     @        i       j                 �|�:@�q�q�?             @        ������������������������       �                      @       ������������������������       �                     �?        ������������������������       �                     @       ������������������������       �                     @        n       o                 ���4@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        q       �                 ��D:@\���(\�?�             y@       r       �                    �?\2R}�?�            r@        s       ~                 �|Y=@�θV�?,            @Q@        t       }                    �?����X�?
             ,@       u       z                    �?�q�q�?             (@       v       w                   �8@�z�G��?             $@        ������������������������       �                     @       x       y                   @@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        {       |                    ;@      �?              @        ������������������������       �                     �?       ������������������������       �                     �?       ������������������������       �                      @              �                 �|�=@�1�`jg�?"            �K@       �       �                    �?Du9iH��?            �E@        �       �                    �?$�q-�?
             *@�z�  ������������������������       �        	             (@ �z�  ������������������������       �                     �?0�}�  �       �                   `3@��S�ۿ?             >@��|�  �       �                 ���@h�����?             <@ �4�  ������������������������       �                     $@ -b}�  �       �                   @'@�X�<ݺ?
             2@�b}�  ������������������������       �$�q-�?             *@p�z�  ������������������������       �                     @p�z�  �       �                    �?      �?              @ p.}�  ������������������������       �                     �?�-z�  ������������������������       �                     �?p�z�  ������������������������       �                     (@i�y�  �       �                   @4@�2�~w�?�            �k@ �z�  �       �                 pf� @      �?             0@ �b}�  �       �                    �?      �?              @?"}�  ������������������������       �                     @��b}�  ������������������������       �                     @ �z�  ������������������������       �                      @�)b}�  �       �                   �<@ =[y��?y            �i@ �3�  ������������������������       �        '            @P@p�z�  �       �                   �*@��X�-�?R            `a@�z�  �       �                     @�#-���?@            @Z@ �3�  �       �                   �F@r�q��?             8@=�y�  �       �                   @D@���y4F�?             3@*b}�  �       �                 `fF)@r�q��?             2@�G}�  ������������������������       �                     $@pw�|�  �       �                 �|�=@      �?              @ �3�  ������������������������       �                      @�z�  �       �                    @@r�q��?             @ w�y�  ������������������������       �                     @��b}�  �       �                   @B@�q�q�?             @�z�  ������������������������       �      �?              @ؼ�  ������������������������       �                     �? �-}�  ������������������������       �                     �?p�z�  ������������������������       �                     @ �b}�  �       �                 ���"@xdQ�m��?/            @T@�.}�  �       �                 ��@ �\���?-            �S@ Zz�  ������������������������       �                     7@plz�  �       �                 ��L@@4և���?!             L@ (z�  �       �                 �|Y>@���Q��?             @ �>~�  ������������������������       �                      @p?z�  ������������������������       �                     @ �z�  �       �                   �@@`'�J�?            �I@I�z�  �       �                 ��) @`Jj��?             ?@�b}�  �       �                 @3�@h�����?             <@lz�  �       �                 �?�@��S�ۿ?             .@�b}�  ������������������������       �                     $@ �b}�  ������������������������       �z�G�z�?             @ �b}�  ������������������������       �                     *@0�z�  �       �                 �|Y=@�q�q�?             @ ��y�  ������������������������       �                     �?0�b}�  �       �                 �|�>@      �?              @ 5�  ������������������������       �                     �?�z�  ������������������������       �                     �?pB7�  ������������������������       �        	             4@p�z�  �       �                    ?@      �?              @ �z�  ������������������������       �                     �?`�b}�  ������������������������       �                     �? Sz�  ������������������������       �                     A@0(z�  �       �                 p�w@�/e�U��?A            �[@�}�  �       �                    �?� �W�??            �Z@�}�  �       �                    �?X�Cc�?4             U@ �z�  �       �                 @�pX@
;&����?             7@�}�  �       �                    �?b�2�tk�?             2@�}�  �       �                 �|�;@�eP*L��?             &@ @/}�  ������������������������       �                      @��:}�  �       �                 ��2>@�q�q�?             "@ �z�  ������������������������       �                      @ �:}�  �       �                    C@؇���X�?             @��  ������������������������       �                     @        �       �                 �D D@�q�q�?             @    n   ������������������������       �                     �?   f   ������������������������       �                      @i   n   �       �                 ��`E@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @v   e   ������������������������       �                     @
       �       �                    R@�ɞ`s�?%            �N@   )   �       �                 03k:@�c�Α�?$             M@    s   ������������������������       �                      @       �       �                 �!fK@      �?#             L@   e   �       �                     �?z�G�z�?             D@   n   �       �                    <@��G���?            �B@    d   ������������������������       �                     �?    f   �       �                   �F@r�q��?             B@   _   �       �                    �?�E��ӭ�?             2@   e   �       �                   `@@�n_Y�K�?
             *@    0   �       �                 �|Y=@r�q��?             @    e   ������������������������       �                     �?a   s   ������������������������       �                     @   "   ������������������������       �                     @u   r   ������������������������       �                     @i   n   �       �                   @J@�X�<ݺ?
             2@    e   �       �                 `f�;@      �?              @    [   ������������������������       �                     �?
       ������������������������       �                     @    n   ������������������������       �                     $@    ,   ������������������������       �                     @_   l   �       �                    �?     ��?             0@   c   �       �                     @�n_Y�K�?	             *@       �       �                    C@�<ݚ�?             "@   t   �       �                 �|Y>@���Q��?             @   b   ������������������������       �                     @    t   ������������������������       �                      @    o   ������������������������       �                     @    m   �       �                    >@      �?             @   d   �       �                    ;@      �?              @    d   ������������������������       �                     �?        ������������������������       �                     �?    a   ������������������������       �                      @    k   �       �                 ���[@�q�q�?             @    '   ������������������������       �                     �?        ������������������������       �                      @l   f   ������������������������       �                     @
       �       �                     �?�nkK�?             7@       �       �                    �?�8��8��?             (@    f   �       �                 ��UO@؇���X�?             @        ������������������������       �                     @   f   �       �                   @D@�q�q�?             @        ������������������������       �                     �?t       ������������������������       �                      @        ������������������������       �                     @i   f   ������������������������       �                     &@   n   ������������������������       �                     @       �t�b�     h�h*h-K ��h/��R�(KK�KK��h]�B�       p{@      q@     �M@     �R@     �A@     @R@      @     �E@              2@      @      9@              2@      @      @              @      @      @      �?      @              @      �?               @              @@      >@      ,@              2@      >@       @              0@      >@      (@      0@      (@      (@      @      @       @              �?      @              @      �?              "@      "@      �?      "@      �?      @              @       @                      @      @      ,@       @               @      ,@              $@       @      @       @      @       @       @       @                       @              �?              �?      8@       @               @      8@             �w@     �h@     �A@     �a@      @     �Y@      @     �X@              A@      @      P@      @     �C@              =@      @      $@      �?               @      $@              @       @      @              @       @                      9@       @      @       @                      @      >@     �C@      9@      C@      6@      C@       @      6@       @      3@       @      $@              �?       @      "@      @       @      @       @               @      @              @              �?      @      �?                      @              "@              @      ,@      0@      &@      0@      $@      $@      @      @      @       @               @      @              �?      @      �?                      @      @      @       @               @      @      �?      @      �?      �?      �?                      �?               @      �?              �?      @              @      �?       @               @      �?              @              @              @      �?              �?      @             �u@     �K@     �p@      4@      O@      @      $@      @       @      @      @      @      @              �?      @      �?                      @      �?      �?      �?                      �?       @              J@      @      D@      @      (@      �?      (@                      �?      <@       @      ;@      �?      $@              1@      �?      (@      �?      @              �?      �?      �?                      �?      (@             �i@      *@      (@      @      @      @      @                      @       @             `h@      "@     @P@             @`@      "@      X@      "@      4@      @      .@      @      .@      @      $@              @      @               @      @      �?      @               @      �?      �?      �?      �?                      �?      @              S@      @     �R@      @      7@              J@      @      @       @               @      @             �H@       @      =@       @      ;@      �?      ,@      �?      $@              @      �?      *@               @      �?      �?              �?      �?              �?      �?              4@              �?      �?              �?      �?              A@              S@     �A@      S@      ?@      K@      >@      (@      &@      @      &@      @      @               @      @      @               @      @      �?      @               @      �?              �?       @              �?      @      �?                      @      @              E@      3@      E@      0@               @      E@      ,@     �@@      @      >@      @              �?      >@      @      *@      @       @      @      �?      @      �?                      @      @              @              1@      �?      @      �?              �?      @              $@              @              "@      @       @      @      @       @      @       @      @                       @      @              �?      @      �?      �?              �?      �?                       @      �?       @      �?                       @              @      6@      �?      &@      �?      @      �?      @               @      �?              �?       @              @              &@                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJW:+LhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM)huh*h-K ��h/��R�(KM)��h|�B@J         r                    �?]@f�
�?�           8�@               a                    �?��K�"�?�            �q@ o u r        &                 `f�$@�e�U��?�            �m@      @       %                    �?��H�}�?              I@              "                    �?(���@��?            �G@     0@                        �̌@���� �?            �D@     @                        ���@�r����?             >@      "@       	                 �|Y:@����X�?             @      @������������������������       �                     @        
                           �?�q�q�?             @        ������������������������       �                     �?       @������������������������       �                      @      @                           �?���}<S�?             7@       ������������������������       �        	             0@      $@                           4@����X�?             @      "@������������������������       �                     �?       @                        �&B@r�q��?             @     C@                          �7@�q�q�?             @      �?������������������������       �                      @       @������������������������       �                     �?        ������������������������       �                     @      0@                          �2@���|���?             &@       @������������������������       �                     �?                                ��� @�z�G��?             $@     @                        @3�@r�q��?             @     �?                          �8@�q�q�?             @      @������������������������       �                     �?                                   ;@      �?              @        ������������������������       �                     �?      @������������������������       �                     �?      @������������������������       �                     @                !                  SE"@      �?             @      @������������������������       �                      @ ���  ������������������������       �                      @�8��  #       $                   �3@�q�q�?             @ ���  ������������������������       �                      @���  ������������������������       �                     @���  ������������������������       �                     @ >��  '       `                 �QD@X�E)9�?v            �g@��  (       E                    �?�<�}���?K            @^@��  )       D                    @�? Da�?(            �O@��  *       +                    �?\#r��?&            �N@ ��  ������������������������       �                     @ ��  ,       5                 `f�)@ �Cc}�?#             L@ ���  -       .                 pF%@`2U0*��?             9@      �?������������������������       �                     *@���  /       0                    +@�8��8��?             (@ ��  ������������������������       �                     @ ���  1       4                    �?r�q��?             @N��  2       3                 ��&@z�G�z�?             @ ���  ������������������������       �                     �?     @������������������������       �                     @���  ������������������������       �                     �?���  6       =                   �*@�חF�P�?             ?@ ���  7       <                   �B@X�<ݚ�?             "@���  8       ;                    �?����X�?             @��  9       :                    <@�q�q�?             @ ���  ������������������������       �                      @ ���  ������������������������       �                     @0��  ������������������������       �                     �? <��  ������������������������       �                      @���  >       ?                    �?���7�?             6@���  ������������������������       �                     .@b��  @       C                    1@؇���X�?             @��  A       B                    "@�q�q�?             @       ������������������������       �                      @      @������������������������       �                     �?     @������������������������       �                     @        ������������������������       �                      @       F       _                   �@@V�a�� �?#             M@       G       H                    �?F�t�K��?"            �L@        ������������������������       �        	             .@       I       J                   �9@0,Tg��?             E@        ������������������������       �                     ,@       K       T                     @��>4և�?             <@       L       M                    6@      �?             0@        ������������������������       �                      @        N       S                    :@؇���X�?
             ,@       O       P                   �8@�<ݚ�?             "@        ������������������������       �                     �?        Q       R                   �E@      �?              @       ������������������������       �                     @       ������������������������       �                      @        ������������������������       �                     @       U       ^                 �̤=@�q�q�?             (@       V       ]                 `fV6@�z�G��?             $@       W       X                 �|�;@և���X�?             @        ������������������������       �                     @        Y       Z                 03�1@      �?             @        ������������������������       �                      @        [       \                 03C3@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?       ������������������������       �        +             Q@       b       q                    @v�2t5�?            �D@       c       d                    �?      �?             A@        ������������������������       �                     @        e       f                     @�f7�z�?             =@        ������������������������       �                     @        g       h                    @�q�q�?             8@        ������������������������       �                     @        i       n                    *@p�ݯ��?
             3@       j       k                    @�8��8��?             (@        ������������������������       �                     @        l       m                    @r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        o       p                 ���4@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?       ������������������������       �                     @        s       �                 ��D:@���<��?           �z@       t       y                    $@�%�P��?�            �t@        u       v                     @"pc�
�?             &@        ������������������������       �                     @        w       x                 ��|2@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        z       �                     @ E�+0+�?�            �s@        {       |                   �)@�(\����?1             T@        ������������������������       �                    �A@       }       �                 ��,@`Ӹ����?            �F@       ~                        �|�<@$�q-�?             :@        ������������������������       �                     ,@       �       �                 �|�=@r�q��?             (@        ������������������������       �                     �?�z�  �       �                   �A@�C��2(�?             &@�z�  �       �                    @@r�q��?             @ �}�  ������������������������       �                      @���|�  ������������������������       �      �?             @ �4�  ������������������������       �                     @0-b}�  ������������������������       �                     3@��b}�  �       �                    �?��5Վ3�?�            �m@ �z�  �       �                    �?^������?            �A@�z�  �       �                    �?�c�Α�?             =@p.}�  �       �                 ���@      �?             8@ -z�  ������������������������       �                     @p�z�  �       �                   @@�q�q�?
             2@ i�y�  �       �                   �5@X�<ݚ�?             "@ �z�  ������������������������       �                      @0�b}�  �       �                 �|=@և���X�?             @ ?"}�  ������������������������       �                      @ �b}�  ������������������������       ����Q��?             @p�z�  �       �                 �|�;@�����H�?             "@ )b}�  �       �                   �2@      �?             @ �3�  ������������������������       �                     @p�z�  ������������������������       �                     �?��z�  ������������������������       �                     @ �3�  �       �                 �&�)@���Q��?             @ =�y�  ������������������������       �                      @*b}�  ������������������������       �                     @�G}�  �       �                 ��y&@�q�q�?             @ w�|�  ������������������������       �                      @0�3�  ������������������������       �                     @p�z�  �       �                   @@@ ��fί�?�            `i@w�y�  �       �                    �?3��e��?j            �d@�b}�  �       �                   �:@$s��O�?Z            �a@ �z�  �       �                   �2@�FVQ&�?,            �P@ ��  �       �                   �1@      �?
             (@�-}�  �       �                   �0@�<ݚ�?             "@�z�  �       �                 pf�@����X�?             @ �b}�  ������������������������       �                      @��.}�  �       �                 pFD!@���Q��?             @ Zz�  ������������������������       ��q�q�?             @ lz�  ������������������������       �                      @ (z�  ������������������������       �                      @�>~�  �       �                 ���@�q�q�?             @ ?z�  ������������������������       �                     �?0�z�  �       �                 ��Y @      �?              @ I�z�  ������������������������       �                     �?�b}�  ������������������������       �                     �? lz�  �       �                    �?@3����?"             K@ �b}�  ������������������������       �                      @аb}�  �       �                 ���@ pƵHP�?!             J@ �b}�  �       �                    7@z�G�z�?             @ �z�  ������������������������       �                      @��y�  �       �                   �8@�q�q�?             @ �b}�  ������������������������       �                     �? 5�  ������������������������       �                      @ �z�  ������������������������       �                    �G@pB7�  �       �                 ��) @��A��?.            �R@�z�  �       �                 @3�@lGts��?$            �K@�z�  �       �                   �>@(L���?            �E@�b}�  �       �                 �|Y=@     ��?             @@ Sz�  �       �                    �?z�G�z�?             @ (z�  ������������������������       �                     �? �}�  ������������������������       �                     @��}�  �       �                 ��(@�>����?             ;@�z�  �       �                 03�@      �?             0@ �}�  ������������������������       �                     @�}�  ������������������������       �"pc�
�?             &@ @/}�  ������������������������       �                     &@��:}�  �       �                   �?@���!pc�?             &@ �z�  �       �                 pff@�q�q�?             @ �:}�  ������������������������       �                     @ ��  ������������������������       �                      @p�b}�  �       �                 �?�@z�G�z�?             @ �b}�  ������������������������       �                      @ �b}�  ������������������������       ��q�q�?             @�a}�  ������������������������       �                     (@p�z�  �       �                 ��)"@p�ݯ��?
             3@ �z�  �       �                 �|Y<@      �?              @ �4�  ������������������������       �                     @0G�z�  �       �                 pf� @�q�q�?             @ �z�  ������������������������       �                     �?�}�  ������������������������       �                      @�`z�  �       �                    �?�C��2(�?             &@ )b}�  ������������������������       �                      @ ܾz�  �       �                    (@�����H�?             "@ �'�  �       �                   �<@z�G�z�?             @ �z�  ������������������������       �                      @p�z�  �       �                 �|Y=@�q�q�?             @ �z�  ������������������������       �                     �? �	z�  ������������������������       �                      @ �	z�  ������������������������       �                     @P�b}�  �       �                    �? 7���B�?             ;@�z�  ������������������������       �                     6@�b}�  �       �                    �?z�G�z�?             @ bz�  ������������������������       �                     �? oz�  ������������������������       �                     @p�z�  ������������������������       �                     B@(z�  �                          �J@*Mp����?J            �Y@��  �       �                 ��";@|jq��?<            �T@ ��  �       �                 03k:@      �?              @ �z�  ������������������������       �                     �?p�z�  �       �                 �|�?@����X�?             @ I7�  ������������������������       �                     �?�G}�  �       �                    �?r�q��?             @ �G}�  ������������������������       �                      @��  �       �                   �C@      �?             @ =�y�  ������������������������       �                     �? ؂z�  �       �                    H@�q�q�?             @=�y�  ������������������������       �      �?              @�=�y�  ������������������������       �                     �? ;�y�  �       �                   �;@L�qA��?5            �R@ w-�  �       �                    6@l��[B��?             =@L7�  �       �                    �?�����?             3@�b}�  ������������������������       �                     "@�z�  �       �                    @���Q��?             $@ N7�  ������������������������       �                     @N7�  �       �                    @�q�q�?             @�y�  �       �                    @���Q��?             @ G}�  ������������������������       �                      @0�y�  ������������������������       �                     @P�'�  ������������������������       �                     �?0i�y�  �       �                    �?ףp=
�?             $@�z�  ������������������������       �                     "@�G}�  ������������������������       �                     �?�Wz�  �                           �?���j��?!             G@O7�  �                         �I@P����?             C@�e�  �                          �?<ݚ)�?             B@�e�  �                         �H@����X�?            �A@�e�                         p�w@     ��?             @@2f�                           �?������?             >@                             `f�B@�GN�z�?             6@                               �A@�eP*L��?	             &@             	                   �?�q�q�?             "@                              �|�=@�q�q�?             @        ������������������������       �                     �?                                �A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        
                        �>@r�q��?             @                               @=@�q�q�?             @        ������������������������       �                     �?                              �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     &@                                 �?      �?              @                             `ށK@և���X�?             @        ������������������������       �                      @                                �G@���Q��?             @                                @C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        !      (                   �?�}�+r��?             3@       "      #                   �?$�q-�?	             *@        ������������������������       �                     @        $      '                 )?@r�q��?             @        %      &                  �Q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h*h-K ��h/��R�(KM)KK��h]�B�       z@     `r@      O@     @k@      C@      i@      2@      @@      .@      @@      &@      >@      @      :@       @      @              @       @      �?              �?       @               @      5@              0@       @      @      �?              �?      @      �?       @               @      �?                      @      @      @              �?      @      @      @      �?       @      �?      �?              �?      �?              �?      �?              @               @       @               @       @              @       @               @      @              @              4@      e@      4@     @Y@       @     �K@      @     �K@              @      @      I@      �?      8@              *@      �?      &@              @      �?      @      �?      @      �?                      @              �?      @      :@      @      @       @      @       @      @       @                      @              �?       @              �?      5@              .@      �?      @      �?       @               @      �?                      @       @              (@      G@      &@      G@              .@      &@      ?@              ,@      &@      1@      @      (@       @               @      (@       @      @              �?       @      @              @       @                      @      @      @      @      @      @      @      @              �?      @               @      �?      �?      �?                      �?      @                       @      �?                      Q@      8@      1@      1@      1@              @      1@      (@              @      1@      @      @              (@      @      &@      �?      @              @      �?              �?      @              �?      @              @      �?              @             0v@      S@      r@     �D@       @      "@              @       @      @              @       @             �q@      @@     �S@       @     �A@             �E@       @      8@       @      ,@              $@       @              �?      $@      �?      @      �?       @              @      �?      @              3@              j@      >@      7@      (@      5@       @      2@      @      @              (@      @      @      @               @      @      @       @               @      @       @      �?      @      �?      @                      �?      @              @       @               @      @               @      @       @                      @      g@      2@     �b@      2@     �^@      1@      O@      @      "@      @      @       @      @       @       @              @       @      �?       @       @               @               @      �?      �?              �?      �?              �?      �?             �J@      �?       @             �I@      �?      @      �?       @               @      �?              �?       @             �G@             �N@      *@     �H@      @     �B@      @      =@      @      @      �?              �?      @              9@       @      ,@       @      @              "@       @      &@               @      @      @       @      @                       @      @      �?       @               @      �?      (@              (@      @       @      @              @       @      �?              �?       @              $@      �?       @               @      �?      @      �?       @               @      �?              �?       @              @              :@      �?      6@              @      �?              �?      @              B@             �P@     �A@     �H@      A@       @      @              �?       @      @      �?              �?      @               @      �?      @              �?      �?       @      �?      �?              �?     �G@      <@      ,@      .@      *@      @      "@              @      @              @      @       @      @       @               @      @              �?              �?      "@              "@      �?             �@@      *@      9@      *@      9@      &@      9@      $@      6@      $@      6@       @      1@      @      @      @      @      @      �?       @              �?      �?      �?      �?                      �?      @      �?       @      �?      �?              �?      �?      �?                      �?      @                       @      &@              @      @      @      @       @               @      @       @      �?              �?       @                       @      �?                       @      @                      �?               @       @              2@      �?      (@      �?      @              @      �?      �?      �?      �?                      �?      @              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJF<KdhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM'huh*h-K ��h/��R�(KM'��h|�B�I                             @	dm#��?�           8�@                                   @     ��?              H@ o u r                         �-]@(;L]n�?             >@     (@������������������������       �                     <@       @                        �(\�?      �?              @        ������������������������       �                     �?      @������������������������       �                     �?      �?       	                    �?�<ݚ�?
             2@       @������������������������       �                     $@       
                        ��T?@      �?              @        ������������������������       �                      @      4@                           @�q�q�?             @     @������������������������       �                     @      ,@������������������������       �                      @              "                  @L@^ɼ���?�           ��@     �?       W                    �?@\L5�T�?�           ؃@      �?       4                     @l��TO��?H            @_@     �?                           �?�M���?(             Q@     �`@                        03�=@�X�<ݺ?             B@      *@                            �?      �?              @      @������������������������       �                      @      �?������������������������       �                     @        ������������������������       �                     <@      �?       )                 �D�G@     ��?             @@     @                          �;@��.k���?             1@      �?������������������������       �                     �?      G@       (                     �?     ��?
             0@     @       '                    �?��
ц��?             *@     *@       &                    C@�q�q�?             (@     @       %                   �A@�eP*L��?             &@     @       $                 ��2>@���Q��?             $@     8@        #                 �ܵ<@      �?              @     @!       "                 X�,@@      �?             @      @������������������������       �                      @      @������������������������       �                      @      @������������������������       �                     @      7@������������������������       �                      @      @������������������������       �                     �?      @������������������������       �                     �?      .@������������������������       �                     �?      @������������������������       �                     @      �?*       +                  �}S@������?
             .@      �?������������������������       �                     @      (@,       3                    �?      �?              @      @-       2                    �?�q�q�?             @     @.       1                    �?      �?             @       /       0                   �=@�q�q�?             @      @������������������������       �                     �?      �?������������������������       �                      @       @������������������������       �                     �?        ������������������������       �                      @       @������������������������       �                      @        5       N                    �?�MWl��?             �L@       6       9                    �?:	��ʵ�?            �F@      �?7       8                 `�@1@      �?              @     K@������������������������       �                     @        ������������������������       �                      @      @:       G                 �|Y=@�MI8d�?            �B@        ;       @                 ���@X�Cc�?             ,@      @<       =                    5@���Q��?             @        ������������������������       �                     �?        >       ?                   �7@      �?             @      �?������������������������       �                     @        ������������������������       �                     �?        A       F                   �<@�<ݚ�?             "@     @B       C                   �8@      �?              @        ������������������������       �                     @        D       E                   @;@�q�q�?             @        ������������������������       �                     �?      @������������������������       �                      @      �?������������������������       �                     �?       @H       I                 ���@�nkK�?             7@        ������������������������       �                     @      �?J       M                 �|�=@      �?             0@       K       L                   @@�C��2(�?             &@       ������������������������       �؇���X�?             @        ������������������������       �                     @        ������������������������       �                     @        O       V                 ���.@�q�q�?             (@       P       U                    �?      �?              @       Q       R                    �?r�q��?             @        ������������������������       �                     @        S       T                 �&�)@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        X                       0�^I@Gq����?F           �@       Y       �                     @�"��c��?           P|@        Z       �                    �?z�7�Z�?\            @b@       [       t                 �|Y=@$��fF?�?L            @_@        \       a                    &@H�z�G�?             D@        ]       ^                    �?X�Cc�?             ,@        ������������������������       �                     @        _       `                   �7@����X�?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        b       k                   �;@�	j*D�?             :@       c       f                    �?�t����?             1@        d       e                    7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        g       h                    :@��S�ۿ?             .@       ������������������������       �        	             (@        i       j                     �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        l       m                    �?�q�q�?             "@        ������������������������       �                     @        n       s                 `f�D@���Q��?             @       o       p                 `fF<@�q�q�?             @        ������������������������       �                     �?        q       r                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        u       �                   �*@ܻ�yX7�?1            @U@        v       }                   �>@��p\�?            �D@        w       x                    �?�r����?
             .@        ������������������������       �                     �?        y       |                 �|�=@@4և���?	             ,@       z       {                    @�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     @        ~                           �? ��WV�?             :@        ������������������������       �                     �?        ������������������������       �                     9@        �       �                   �2@���|���?             F@    )   ������������������������       �                     @ D]i 
 ��       �                   @J@�z�G��?             D@   .   �       �                    �?�q�q�?             B@   t   �       �                    �?`�Q��?             9@        ������������������������       �                      @        �       �                     �?��+7��?             7@   g   �       �                   �>@�z�G��?             4@   "   �       �                 ��<:@�eP*L��?             &@        ������������������������       �                      @   f   �       �                 X��B@�q�q�?             "@    s   ������������������������       �                      @   b   �       �                    H@և���X�?             @       ������������������������       �      �?             @       ������������������������       �                     �?        ������������������������       �                     "@    b   ������������������������       �                     @   _   �       �                    �?���|���?             &@        �       �                   �E@�q�q�?             @       ������������������������       �                     @   t   ������������������������       �                      @       ������������������������       �                     @    =   ������������������������       �                     @   p   �       �                    *@���N8�?             5@    
   ������������������������       �                      @    s   �       �                    �?�S����?             3@   =   ������������������������       �                     0@       ������������������������       �                     @    s   �       �                    �?4����?�            0s@    u   �       �                    �?      �?             L@        �       �                    @���B���?             :@   e   �       �                    �?���}<S�?             7@   s   �       �                 �|�9@      �?	             0@    e   ������������������������       �                     @       �       �                  ��@z�G�z�?             $@    r   ������������������������       �                      @   n   ������������������������       �                      @   s   ������������������������       �                     @        ������������������������       �                     @o   k   ������������������������       �                     >@       �       �                    �?���w;�?�            `o@        �       �                    �?�G�5��?)            @Q@       �       �                 ���1@b�2�tk�?             B@   e   �       �                 �|�<@��S���?             >@   n   �       �                 pf�@�q�q�?             2@    o   ������������������������       �                     @        �       �                   �2@z�G�z�?	             .@        ������������������������       �                     @    l   �       �                    �?      �?             (@   b   �       �                   �@�<ݚ�?             "@    o   �       �                 �&B@�q�q�?             @       �       �                   �7@      �?              @    h   ������������������������       �                     �?    g   ������������������������       �                     �?   w   ������������������������       �                     �?        ������������������������       �                     @    e   �       �                 �!@�q�q�?             @    N   ������������������������       �                     �?o   n   ������������������������       �                      @    t   �       �                    �?�q�q�?	             (@    H   �       �                   &@      �?             @   ,   ������������������������       �                     @    a   ������������������������       �                     �?       �       �                 ��Y.@      �?              @    e   ������������������������       �                     �?       ������������������������       �                     @    r   ������������������������       �                     @   P   �       �                    :@�C��2(�?            �@@       �       �                   �6@@�0�!��?
             1@   k   �       �                   �0@��S�ۿ?	             .@   e   ������������������������       �                     "@   e   �       �                    3@r�q��?             @    a   ������������������������       �                     �?    c   ������������������������       �                     @    e   ������������������������       �                      @    a   ������������������������       �                     0@        �       �                 �?�@|)����?z            �f@    a   �       �                    ?@@�)�n�?9            @U@   n   �       �                    �?�\=lf�?-            �P@   v   �       �                 ���@ ������?)            �O@    a   �       �                   �8@�����H�?             "@    c   �       �                   �4@z�G�z�?             @    s   ������������������������       �                     �?   i   �       �                 �&b@      �?             @    e   ������������������������       �                     @    x   ������������������������       �                     �?       ������������������������       �                     @   n   ������������������������       �        #             K@   l   ������������������������       �                     @        �       �                 �&B@�����H�?             2@   a   ������������������������       �                     (@       �       �                   �A@�q�q�?             @        �       �                   �@      �?             @    h   ������������������������       �                      @   a   ������������������������       �                      @        ������������������������       �                      @   e   �                          �?�*v��?A            @X@       �       �                 @3�@ ��~���?<            �V@    I   �       �                    �?X�Cc�?             ,@       �       �                   �A@�	j*D�?             *@       �       �                   �:@"pc�
�?             &@    c   ������������������������       �                     @    a   ������������������������       ����Q��?             @    f   ������������������������       �                      @        ������������������������       �                     �?   e   �       �                    )@�KM�]�?4             S@    o   ������������������������       �                     �?   "   �                          ?@���Lͩ�?3            �R@   o   �                       �|�=@H�ՠ&��?$             K@   ,   �                          �?���C��?#            �J@       �                          �?�t����?!            �I@   e   �                       @3�!@(L���?            �E@   E   �       �                 �|Y<@@�0�!��?             A@   _   �       �                 pf� @      �?             0@   e   �       �                 0S5 @"pc�
�?	             &@   x   �       �                   �3@�<ݚ�?             "@    ,   �       �                   �1@      �?             @    h   ������������������������       �                     �?    
   ������������������������       ��q�q�?             @        ������������������������       �                     @   o   ������������������������       �                      @    t   �       �                    8@���Q��?             @   t   ������������������������       �                     @"   
   ������������������������       �                      @    t   �       �                 ��) @�����H�?
             2@       ������������������������       �                     .@    ,   �                        pf� @�q�q�?             @    s   ������������������������       �                      @       ������������������������       �                     �?       ������������������������       �                     "@       ������������������������       �                      @       ������������������������       �                      @       ������������������������       �                     �?       ������������������������       �                     5@       ������������������������       �                     @                                 @�q�q�?*            �L@       	      
                   �?���3�E�?%             J@       ������������������������       �                     @@                                �?      �?             4@Z _b��                           �?�E��ӭ�?             2@                               �E@     ��?             0@                              x#J@�n_Y�K�?             *@        ������������������������       �                     @                                 �?      �?             $@        ������������������������       �                     �?                              `�iJ@X�<ݚ�?             "@        ������������������������       �                     @                              `f�N@�q�q�?             @                                7@      �?             @        ������������������������       �                     �?                                 A@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @              !                   �?z�G�z�?             @                                  ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        #      &                   �?h�����?             <@        $      %                  pE@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     :@        �t�bh�h*h-K ��h/��R�(KM'KK��h]�Bp       0}@     �n@      .@     �@@      �?      =@              <@      �?      �?              �?      �?              ,@      @      $@              @      @       @               @      @              @       @             @|@     `j@     �z@     @j@     �M@     �P@      .@     �J@       @      A@       @      @       @                      @              <@      *@      3@      "@       @              �?      "@      @      @      @      @      @      @      @      @      @       @      @       @       @       @                       @              @       @              �?                      �?      �?              @              @      &@              @      @      @      @       @       @       @      �?       @      �?                       @      �?               @                       @      F@      *@     �B@       @      @       @      @                       @      ?@      @      "@      @       @      @      �?              �?      @              @      �?              @       @      @      �?      @               @      �?              �?       @                      �?      6@      �?      @              .@      �?      $@      �?      @      �?      @              @              @      @      @      �?      @      �?      @              �?      �?              �?      �?               @                      @     �v@      b@     �u@     �Z@     �W@      J@     @V@      B@      7@      1@      @      "@              @      @       @      �?       @      @              2@       @      .@       @      �?      �?              �?      �?              ,@      �?      (@               @      �?              �?       @              @      @              @      @       @      �?       @              �?      �?      �?              �?      �?               @             �P@      3@      C@      @      *@       @              �?      *@      �?      $@      �?      $@                      �?      @              9@      �?              �?      9@              <@      0@              @      <@      (@      8@      (@      1@       @               @      1@      @      ,@      @      @      @       @              @      @               @      @      @      @      @              �?      "@              @              @      @       @      @              @       @              @              @              @      0@       @              @      0@              0@      @             �o@      K@     �A@      5@      @      5@       @      5@       @      ,@              @       @       @       @                       @              @      @              >@             @k@     �@@      J@      1@      6@      ,@      0@      ,@      (@      @              @      (@      @      @              "@      @      @       @      �?       @      �?      �?              �?      �?                      �?      @               @      �?              �?       @              @       @      @      �?      @                      �?      �?      @      �?                      @      @              >@      @      ,@      @      ,@      �?      "@              @      �?              �?      @                       @      0@             �d@      0@     �T@      @     �P@      �?      O@      �?       @      �?      @      �?      �?              @      �?      @                      �?      @              K@              @              0@       @      (@              @       @       @       @               @       @               @              U@      *@     @S@      *@      "@      @      "@      @      "@       @      @              @       @               @              �?      Q@       @              �?      Q@      @     �G@      @     �G@      @     �F@      @     �B@      @      <@      @      (@      @      "@       @      @       @       @       @      �?              �?       @      @               @              @       @      @                       @      0@       @      .@              �?       @               @      �?              "@               @               @                      �?      5@              @              3@      C@      .@     �B@              @@      .@      @      *@      @      &@      @       @      @      @              @      @      �?              @      @              @      @       @       @       @      �?              �?       @               @      �?               @              @               @               @              @      �?      �?      �?              �?      �?              @              ;@      �?      �?      �?      �?                      �?      :@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJؽ�hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B�C         P                     �?e�L��?�           8�@     �F@       3                    �?�G�z�?f             d@ o u r                            �?���r
��?A            @X@ y��                             �?�D����?             E@   p y                           @H@p�ݯ��?             C@     @                        �|�;@�������?             >@      3@������������������������       �                     &@      @       	                    �?p�ݯ��?             3@     @������������������������       �                     $@        
                          �A@�<ݚ�?             "@                               X�,@@����X�?             @                               ��2>@r�q��?             @      @������������������������       �                     �?      @������������������������       �                     @      �?������������������������       �                     �?        ������������������������       �                      @      �?                        ��Z@      �?              @     �?������������������������       �                     @      @������������������������       �                     �?      @                        �\@      �?             @      �?������������������������       �                     �?      �?������������������������       �                     @      �?       *                 0�_J@N{�T6�?$            �K@                                  �?��.k���?             A@        ������������������������       �                     @                               �|�<@���Q��?             >@      @������������������������       �                     @      @       )                    R@�q�q�?             ;@      @       (                    L@�	j*D�?             :@              '                   �>@���Q��?             4@      @                         �̌*@�q�q�?             (@      >@������������������������       �                      @      @!       "                   �C@z�G�z�?             $@      (@������������������������       �                     @      @#       &                 `f�;@�q�q�?             @      @$       %                    H@z�G�z�?             @       ������������������������       �      �?             @      @������������������������       �                     �?      0@������������������������       �                     �?        ������������������������       �                      @      5@������������������������       �                     @        ������������������������       �                     �?        +       0                 03c@؇���X�?             5@     ,@,       -                    �?�IєX�?	             1@       ������������������������       �                     .@      �?.       /                    =@      �?              @        ������������������������       �                     �?       @������������������������       �                     �?      @1       2                 ���f@      �?             @      @������������������������       �                      @      �?������������������������       �                      @        4       O                   �P@�<ݚ�?%            �O@     �?5       @                 ��Q@���*�?$             N@      �?6       7                    �?�q�q�?             2@        ������������������������       �                     @       @8       ?                    F@�eP*L��?             &@       9       :                    �?r�q��?             @      @������������������������       �                      @       @;       >                   @B@      �?             @     @<       =                   @K@�q�q�?             @      @������������������������       �                     �?       @������������������������       �                      @        ������������������������       �                     �?       @������������������������       �                     @       @A       H                    �?���H��?             E@     @B       G                    �?`Jj��?             ?@     @C       D                    �?$�q-�?             :@       ������������������������       �        
             2@      @E       F                 ���^@      �?              @     �?������������������������       �                     @       @������������������������       �                      @        ������������������������       �                     @      @I       L                    �?���!pc�?             &@       J       K                 �U�X@؇���X�?             @     �?������������������������       �                     @       @������������������������       �                     �?      �?M       N                 ��f`@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        Q       �                    �?�w�+`�?]           8�@       R       �                 Ь�#@�;�T<:�?           �z@       S       T                 ���@D�a�ў�?�            �p@        ������������������������       �                     <@        U       V                 ��@�.�PI�?�            �m@        ������������������������       �                     @        W       X                    /@P�z�?�            `m@        ������������������������       �                      @        Y       p                    �?F�|���?�             m@        Z       [                    �?Dc}h��?&             L@        ������������������������       �        	             *@        \       i                    �?�ʈD��?            �E@       ]       h                 �� @�LQ�1	�?             7@       ^       a                 ���@؇���X�?             5@        _       `                 �|�9@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        b       g                 �|Y=@r�q��?	             (@        c       d                   @8@�q�q�?             @        ������������������������       �                     �?        e       f                   @@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @        j       k                 ���@P���Q�?             4@        ������������������������       �                     @        l       o                 X�I@      �?             0@       m       n                 ��(@��S�ۿ?             .@       ������������������������       �$�q-�?             *@        ������������������������       �                      @        ������������������������       �                     �?        q       v                    �?$���?f             f@        r       u                   �@
;&����?             7@        s       t                   �A@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                     &@        w       �                 �?�@�C��2(�?Z            @c@       x       y                 �|�<@����D��?5            @W@       ������������������������       �                     J@        z       �                   @@@������?            �D@       {       �                   �@�8��8��?             8@        |       �                 �&B@����X�?             @       }       ~                 ��@r�q��?             @        ������������������������       �                     @               �                 �|Y>@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?       ������������������������       �                     �?    p   ������������������������       �        	             1@    s   ������������������������       �                     1@    f   �       �                   �4@`��:�?%            �N@        �       �                   �0@�q�q�?
             .@        ������������������������       ����Q��?             @        �       �                 @3�@�z�G��?             $@    n   ������������������������       �                      @        �       �                 ��Y @      �?              @    o   �       �                   �2@      �?             @    t   ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @   s   �       �                 @3�@*
;&���?             G@    S   �       �                   �A@      �?              @        ������������������������       �      �?             @   T   ������������������������       �      �?              @   t   �       �                    �?�˹�m��?             C@   y   �       �                 �|Y=@�8��8��?             B@    t   ������������������������       �                     "@        �       �                 �|Y?@�����H�?             ;@   ,   �       �                 ��) @r�q��?	             2@   y   ������������������������       �                     &@        �       �                 pf� @և���X�?             @    o   ������������������������       �                     @       ������������������������       �                     @    n   ������������������������       �                     "@   m   ������������������������       �                      @    i   �       �                   �F@v�_���?e            �c@       �       �                   P,@�S��<�?Y            �a@    e   �       �                    �?      �?$             N@    
   �       �                     @ 7���B�?             ;@       ������������������������       �                     4@   _   �       �                    �?؇���X�?             @       �       �                 �[$@r�q��?             @        ������������������������       �                     @    i   �       �                 ��&@�q�q�?             @    y   ������������������������       �                     �?        ������������������������       �                      @    n   ������������������������       �                     �?   o   �       �                 �%@<���D�?            �@@    b   ������������������������       �                     @       �       �                     @8�Z$���?             :@       �       �                 �|�<@�8��8��?             8@   t   ������������������������       �                     &@       �       �                 �|�=@8�Z$���?             *@        ������������������������       �                      @   l   ������������������������       �                     &@   .   ������������������������       �                      @    n   �       �                 pf�/@d�� z�?5            @T@        �       �                    1@      �?             0@        �       �                   �-@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?    v   ������������������������       �        
             ,@       �       �                     @�4��?)            @P@       �       �                    �?؀�:M�?            �B@        �       �                    �?      �?
             0@    e   ������������������������       �                     @    a   �       �                    �?z�G�z�?             $@        ������������������������       �                     @    v   �       �                   �;@����X�?             @        ������������������������       �                     �?       �       �                   �E@r�q��?             @   F   ������������������������       �                     @       ������������������������       �                     �? K@lt �������������������������       �                     5@    
   �       �                 ���1@����X�?             <@        �       �                    �?      �?              @   ,   ������������������������       �                     @G   r   ������������������������       �                     @       �       �                    �?R���Q�?             4@    r   �       �                   �2@      �?              @    t   ������������������������       �                     @   c   �       �                    �?���Q��?             @        ������������������������       �                      @    i   �       �                 �|�;@�q�q�?             @    p   ������������������������       �                     �?    )   ������������������������       �                      @       ������������������������       �                     (@    l   �       �                   �.@�IєX�?             1@       ������������������������       �        	             ,@   t   �       �                    5@�q�q�?             @    a   ������������������������       �                     �?        ������������������������       �                      @   p   �       �                     @X9����?U            �_@        �       �                   �6@�������?             A@        ������������������������       �        
             .@   t   �       �                 ��J@�\��N��?             3@   e   �       �                    @���Q��?             .@       �       �                    �?X�Cc�?             ,@        ������������������������       �                     @       ������������������������       �                     "@        ������������������������       �                     �?       ������������������������       �                     @   t   �       �                    �?R�(��?=            @W@        �       �                 X��B@���y4F�?             3@       �       �                    @r�q��?             2@       �       �                    �?d}h���?             ,@       �       �                    3@r�q��?	             (@   e   �       �                    &@�q�q�?             @   n   ������������������������       �                     @    x   ������������������������       �                      @    i   ������������������������       �                     @       �       �                 �|Y=@      �?              @    #   ������������������������       �                     �?    .   ������������������������       �                     �?    t   ������������������������       �                     @    t   ������������������������       �                     �?       �                       �̼6@^��4m�?0            �R@        �                       �̌5@�'�=z��?            �@@   a   �       �                   �*@*;L]n�?             >@    r   �       �                    (@�z�G��?             $@       ������������������������       �                     @       �       �                 xFT$@���Q��?             @        ������������������������       �                     @   _   ������������������������       �                      @       �       �                    �?�z�G��?             4@       �       �                     @8�Z$���?	             *@       �       �                    )@"pc�
�?             &@        ������������������������       �                      @    s   ������������������������       �                     "@    a   ������������������������       �                      @   r   �       �                 @33/@և���X�?             @        ������������������������       �                     �?        �                           �?�q�q�?             @        ������������������������       �                     @                                 +@�q�q�?             @        ������������������������       �                     �?       ������������������������       �                      @       ������������������������       �                     @             
                   �?��p\�?            �D@              	                  @C@�t����?
             1@                                �B@      �?              @       ������������������������       �                     @       ������������������������       �                      @       ������������������������       �                     "@                             ��p@@ �q�q�?             8@ U =b��                       ��T?@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �        
             *@        �t�b��     h�h*h-K ��h/��R�(KMKK��h]�B�       �{@     �p@      J@      [@      C@     �M@      1@      9@      ,@      8@      @      7@              &@      @      (@              $@      @       @      @       @      @      �?              �?      @                      �?       @              @      �?      @                      �?      @      �?              �?      @              5@      A@      2@      0@              @      2@      (@              @      2@      "@      2@       @      (@       @      @       @       @               @       @              @       @      @      �?      @      �?      @              �?      �?               @              @                      �?      @      2@      �?      0@              .@      �?      �?              �?      �?               @       @       @                       @      ,@     �H@      &@     �H@      @      (@              @      @      @      �?      @               @      �?      @      �?       @      �?                       @              �?      @              @     �B@       @      =@       @      8@              2@       @      @              @       @                      @      @       @      �?      @              @      �?               @       @       @                       @      @             px@      d@     0t@     @Y@     `k@     �G@      <@             �g@     �G@              @     �g@      F@               @     �g@      E@     �C@      1@              *@     �C@      @      4@      @      2@      @       @      �?              �?       @              $@       @      �?       @              �?      �?      �?      �?                      �?      "@               @              3@      �?      @              .@      �?      ,@      �?      (@      �?       @              �?              c@      9@      (@      &@      �?      &@              &@      �?              &@             �a@      ,@     �V@       @      J@             �C@       @      6@       @      @       @      @      �?      @               @      �?      �?      �?      �?                      �?      1@              1@             �H@      (@      $@      @      @       @      @      @               @      @      �?      @      �?              �?      @              @             �C@      @      @      @      @      @      �?      �?     �A@      @     �@@      @      "@              8@      @      .@      @      &@              @      @              @      @              "@               @              Z@      K@      V@     �J@      >@      >@      �?      :@              4@      �?      @      �?      @              @      �?       @      �?                       @              �?      =@      @      @              6@      @      6@       @      &@              &@       @               @      &@                       @      M@      7@      .@      �?      �?      �?      �?                      �?      ,@             �E@      6@      7@      ,@       @      ,@              @       @       @              @       @      @      �?              �?      @              @      �?              5@              4@       @      @      @              @      @              1@      @      @      @      @               @      @               @       @      �?              �?       @              (@              0@      �?      ,@               @      �?              �?       @              Q@     �M@      "@      9@              .@      "@      $@      "@      @      "@      @              @      "@                      �?              @     �M@      A@      @      .@      @      .@      @      &@       @      $@       @      @              @       @                      @      �?      �?              �?      �?                      @      �?             �K@      3@      1@      0@      1@      *@      @      @              @      @       @      @                       @      ,@      @      &@       @      "@       @               @      "@               @              @      @      �?               @      @              @       @      �?              �?       @                      @      C@      @      .@       @      @       @      @                       @      "@              7@      �?      $@      �?      $@                      �?      *@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJX��vhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B@A         d                    �?e�L��?�           8�@               _                    @<�T]���?�            �o@              \                    @Q��"�?�            `m@     @       G                 �|�=@��^���?�             m@     �?                           !@ܱ#_��?\            `b@      �?������������������������       �                     ,@      0@                           '@���c�?T            �`@      "@������������������������       �                     @        	                            @:�����?R            �_@        
                           �?���J��?"            �I@        ������������������������       �                     4@       @                           �?�g�y��?             ?@     @                           9@P���Q�?             4@                                   �?      �?             @     $@                          �'@      �?              @      "@������������������������       �                     �?       @������������������������       �                     �?     �?������������������������       �                      @     �`@������������������������       �                     0@      *@������������������������       �                     &@      @       :                    �?���=A�?0             S@     �?       %                 @� @     ��?)             P@                                 �6@��s����?             E@      �?������������������������       �        
             4@     @                          �9@���|���?             6@      �?                        pf�@      �?             @      G@������������������������       �                     �?     @������������������������       �                     @     *@                           ;@�E��ӭ�?             2@      @������������������������       �                      @     @       $                    �?     ��?             0@     8@        #                 ���@d}h���?	             ,@      @!       "                 �Y�@���Q��?             @        ������������������������       �                      @      >@������������������������       �                     @        ������������������������       �                     "@      @������������������������       �                      @      �?&       1                    �?8�A�0��?             6@       @'       (                   �,@      �?             (@        ������������������������       �                      @      1@)       0                    �?�z�G��?             $@      @*       /                  S�-@�q�q�?             "@       +       .                 �|Y6@���Q��?             @     �?,       -                   �-@�q�q�?             @        ������������������������       �                     �?      �?������������������������       �                      @      *@������������������������       �                      @      �?������������������������       �                     @       @������������������������       �                     �?      @2       9                 �|�:@���Q��?	             $@     �?3       8                    �?؇���X�?             @     @4       5                  �#@      �?             @      �?������������������������       �                      @      �?6       7                 �[$@      �?              @      �?������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @      �?������������������������       �                     @       @;       @                   �6@�q�q�?             (@      �?<       ?                   �3@z�G�z�?             @     @=       >                    �?      �?             @       @������������������������       �                     @        ������������������������       �                     �?      *@������������������������       �                     �?      $@A       B                 �|�:@և���X�?             @      @������������������������       �                      @     @C       D                    �?z�G�z�?             @        ������������������������       �                      @      @E       F                    �?�q�q�?             @      �?������������������������       �                     �?       @������������������������       �                      @        H       W                    �?�̨�`<�?8            @U@     @I       J                   @B@؇���X�?%             L@       ������������������������       �                     ;@     �?K       V                 83'E@�c�Α�?             =@      @L       O                     �?      �?	             0@      �?M       N                    �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        P       U                   �+@�<ݚ�?             "@       Q       T                     @�q�q�?             @       R       S                    D@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     *@        X       Y                     @XB���?             =@       ������������������������       �                     7@        Z       [                    C@r�q��?             @        ������������������������       �                     @        ������������������������       �                     �?       ]       ^                 ��T?@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        `       a                      @�t����?             1@        ������������������������       �                     @        b       c                 �|Y?@$�q-�?
             *@       ������������������������       �        	             (@        ������������������������       �                     �?        e       �                 ��K.@�#2����?"           �|@       f       w                    �?�]l*7��?�            0r@        g       h                   �6@>���Rp�?             M@        ������������������������       �                     "@        i       n                 �|Y=@ i���t�?            �H@        j       m                    �?      �?             (@       k       l                   �<@�q�q�?             "@       ������������������������       �                     @       ������������������������       �                     @       ������������������������       �                     @        o       p                 ���@@-�_ .�?            �B@        ������������������������       �                     .@        q       r                     @�C��2(�?             6@        ������������������������       �                     @        s       v                 �|�=@�����H�?	             2@       t       u                   @@"pc�
�?             &@       ������������������������       �����X�?             @        ������������������������       �                     @        ������������������������       �                     @       x       �                    �?`�q��־?�             m@       y       �                 ���"@ �Cc��?�             l@       z       �                 ��@�1��?o            �e@        {       |                     @��v$���?*            �N@        ������������������������       �                     $@       }       �                 ���@���J��?#            �I@        ~                        ���@�IєX�?
             1@       ������������������������       �        	             0@       ������������������������       �                     �?        ������������������������       �                     A@��z�  �       �                    �?�h����?E             \@Wz�  �       �                   �3@ ѯ��?B            �Z@ ��z�  �       �                   �1@��2(&�?             6@ Xz�  ������������������������       �                     &@TMy� ��       �                 �?�@���!pc�?             &@ �z�  ������������������������       �                     @ �z�  �       �                 ��Y @���Q��?             @Sz�  �       �                   �2@      �?             @ Uz�  ������������������������       �                      @Qz�  ������������������������       �      �?              @ Uz�  ������������������������       �                     �? Vz�  �       �                 �|Y=@@�)�n�?6            @U@ Uz�  ������������������������       �                    �B@ Wz�  �       �                   @@@      �?             H@�z�  �       �                    ?@�#-���?            �A@�z�  �       �                 �|�=@@4և���?             <@�z�  �       �                  sW@HP�s��?             9@ ��z�  ������������������������       �      �?             @�z�  ������������������������       �                     5@ �z�  ������������������������       �                     @ �z�  �       �                 P�@؇���X�?             @ �z�  ������������������������       �                     �?��z�  ������������������������       �                     @ ��z�  ������������������������       �                     *@ �z�  ������������������������       �                     @ �z�  �       �                   @B@�t����?$            �I@�z�  �       �                   �@@R���Q�?             D@l�y�  �       �                     @�ݜ�?            �C@Uz�  �       �                    5@���7�?             6@ Qz�  �       �                   �2@z�G�z�?             @ Wz�  ������������������������       �                      @ �z�  ������������������������       ��q�q�?             @ �z�  ������������������������       �                     1@ �z�  �       �                 `�X#@������?             1@��z�  �       �                   �<@�	j*D�?             *@ �z�  ������������������������       �                     @��z�  �       �                 �|Y=@X�<ݚ�?             "@ �z�  ������������������������       �                      @ Tz�  �       �                 �|�=@����X�?             @ Vz�  ������������������������       �                     @ ��z�  �       �                   �?@      �?             @ ��z�  ������������������������       �                      @ �z�  ������������������������       �                      @ �z�  ������������������������       �                     @ Rz�  ������������������������       �                     �?Uz�  ������������������������       �                     &@ Wz�  �       �                    �?�<ݚ�?             "@ �z�  ������������������������       �                      @ ��z�  �       �                    �?����X�?             @�z�  �       �                     @���Q��?             @ Tz�  ������������������������       �                      @Vz�  ������������������������       �                     @ ��z�  ������������������������       �                      @Uz�  �       �                   �A@      �?l             e@Wz�  �       �                   @A@�Sb(�	�?D             [@j�y�  �       �                 `�/@�Y|���?A            �Y@ ��z�  ������������������������       �                     @ ��z�  �       �                    @�D��??            �X@�z�  �       �                    �?^H���+�?3            �R@Vz�  �       �                    �?�Gi����?            �B@Wz�  �       �                    �?���|���?            �@@ �z�  �       �                      @�q�q�?             "@Qz�  �       �                 �|Y<@����X�?             @ Wz�  �       �                    9@�q�q�?             @ �z�  ������������������������       �                     �? �z�  ������������������������       �                      @�z�  ������������������������       �                     @�z�  �       �                   �2@      �?              @ �z�  ������������������������       �                     �?Uz�  ������������������������       �                     �? l�y�  �       �                   �?@      �?             8@Wz�  �       �                 `f�D@����X�?             5@Wz�  �       �                     �?��
ц��?	             *@Sz�  �       �                   �<@�q�q�?             "@ �z�  ������������������������       �                      @�z�  �       �                 `fF<@և���X�?             @ Wz�  ������������������������       �                      @ �z�  �       �                 �|Y=@z�G�z�?             @ �z�  ������������������������       �                     �?�z�  ������������������������       �                     @�z�  ������������������������       �                     @Tz�  ������������������������       �                      @Vz�  ������������������������       �                     @��z�  �       �                 h"_@      �?             @�z�  ������������������������       �                     @��z�  ������������������������       �                     �?�z�  �       �                    �?V������?            �B@ �z�  �       �                    �?�<ݚ�?             "@��z�  �       �                    ;@      �?              @Wz�  �       �                    �?���Q��?             @�z�  �       �                 8�T@      �?             @ ��z�  ������������������������       �                      @Uz�  ������������������������       �                      @Wz�  ������������������������       �                     �? �z�  ������������������������       �                     @ �z�  ������������������������       �                     �? �z�  �       �                    )@��X��?             <@ m�y�  ������������������������       �                     @ �z�  �       �                 `fFJ@�����?             5@�z�  ������������������������       �        
             .@�z�  �       �                     �?�q�q�?             @�z�  �       �                    7@�q�q�?             @ i�y�  ������������������������       �                     �?    s   ������������������������       �                      @    #   ������������������������       �                     @   k   ������������������������       �                     8@    g   �       �                     �?z�G�z�?             @   i   ������������������������       �                     @    b   ������������������������       �                     �?        �                          �?�?�P�a�?(             N@   p   �       �                    H@r�q��?             E@   t   �       �                    �?`2U0*��?             9@   f   �       �                    �?      �?	             0@    g   ������������������������       �                     �?    _   �       �                   �F@��S�ۿ?             .@    l   �       �                 `fF:@r�q��?             @        ������������������������       �                     @    s   ������������������������       ��q�q�?             @   a   ������������������������       �                     "@       ������������������������       �                     "@   a   �                       �5L@ҳ�wY;�?             1@       �                        i?@������?
             .@       �       �                 `fF:@���|���?             &@    a   ������������������������       �                     @   f   �       �                    �?      �?              @    e   ������������������������       �                     �?                                  L@և���X�?             @    t   ������������������������       �                     @       ������������������������       �                     @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     2@        �t�bh�h*h-K ��h/��R�(KMKK��h]�BP       �{@     �p@     �K@     �h@     �E@      h@     �D@     �g@      @@     �\@              ,@      @@     @Y@      @              :@     @Y@      �?      I@              4@      �?      >@      �?      3@      �?      @      �?      �?              �?      �?                       @              0@              &@      9@     �I@      1@     �G@       @      A@              4@       @      ,@      @      �?              �?      @              @      *@               @      @      &@      @      &@      @       @               @      @                      "@       @              "@      *@      @      "@               @      @      @      @      @      @       @      �?       @      �?                       @       @                      @              �?      @      @      @      �?      @      �?       @              �?      �?              �?      �?              @                      @       @      @      @      �?      @      �?      @                      �?      �?              @      @               @      @      �?       @               @      �?              �?       @              "@      S@       @      H@              ;@       @      5@       @       @      �?      @      �?                      @      @       @      @       @      @       @      @                       @      �?              @                      *@      �?      <@              7@      �?      @              @      �?               @      �?       @                      �?      (@      @              @      (@      �?      (@                      �?     @x@     �Q@     `p@      =@      F@      ,@              "@      F@      @      "@      @      @      @      @                      @      @             �A@       @      .@              4@       @      @              0@       @      "@       @      @       @      @              @             @k@      .@     `j@      *@     �d@      @      N@      �?      $@              I@      �?      0@      �?      0@                      �?      A@             �Z@      @     @Y@      @      3@      @      &@               @      @      @               @      @      �?      @               @      �?      �?      �?             �T@      @     �B@             �F@      @      @@      @      :@       @      7@       @       @       @      5@              @              @      �?              �?      @              *@              @             �F@      @      A@      @      A@      @      5@      �?      @      �?       @               @      �?      1@              *@      @      "@      @      @              @      @               @      @       @      @               @       @               @       @              @                      �?      &@              @       @       @              @       @      @       @               @      @               @             �_@      E@     @R@     �A@      R@      ?@              @      R@      :@      H@      :@      6@      .@      5@      (@      @      @      @       @      �?       @      �?                       @      @              �?      �?      �?                      �?      .@      "@      .@      @      @      @      @      @               @      @      @       @              �?      @      �?                      @      @               @                      @      �?      @              @      �?              :@      &@      @       @      @       @      @       @       @       @               @       @              �?              @              �?              3@      "@              @      3@       @      .@              @       @      �?       @      �?                       @      @              8@              �?      @              @      �?             �J@      @     �A@      @      8@      �?      .@      �?      �?              ,@      �?      @      �?      @               @      �?      "@              "@              &@      @      &@      @      @      @      @              @      @      �?              @      @              @      @              @                       @      2@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ���EhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B�G         r                     @�����?�           8�@                                   �?yÏP�?�            �t@                                03�<@@+K&:~�?[             c@      >@                           �?Xny��?(            �N@     �?                          �H@>A�F<�?             C@     &@                           �?�t����?             A@     4@                          @B@�nkK�?             7@       ������������������������       �                     2@      &@	       
                   �,@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @       @                           �?���!pc�?             &@      @������������������������       �                     �?                                  �;@�z�G��?             $@      $@                          �7@�q�q�?             @      "@������������������������       �                      @       @������������������������       �                     �?     �?                           D@؇���X�?             @     @������������������������       �                     @      @������������������������       �                     �?      �?                           �?      �?             @      �?������������������������       �                      @      �?                          �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?       ������������������������       �                     7@      @������������������������       �        3            �V@      @       =                    �?:���١�?p             f@       @       8                     �?�[�IJ�?            �G@              5                    �?      �?             C@      @                         ��";@��>4և�?             <@      >@������������������������       �                      @      @!       4                 �̾w@$��m��?             :@       "       '                 �|Y<@`�Q��?             9@      >@#       &                    �?      �?              @       $       %                  �}S@և���X�?             @     @������������������������       �                     @      �?������������������������       �                     @       @������������������������       �                     �?        (       3                    �?@�0�!��?             1@     1@)       2                 p�i@@�θ�?	             *@      @*       /                   �A@և���X�?             @       +       ,                 ���<@      �?             @      �?������������������������       �                      @        -       .                 ��2>@      �?              @      �?������������������������       �                     �?      *@������������������������       �                     �?      �?0       1                  �>@�q�q�?             @       @������������������������       �                     �?      @������������������������       �                      @     �?������������������������       �                     @     @������������������������       �                     @      �?������������������������       �                     �?      �?6       7                 ��>Y@z�G�z�?             $@     �?������������������������       �                      @        ������������������������       �                      @        9       :                    �?�����H�?             "@     �?������������������������       �                     @       @;       <                 pV�C@      �?              @      �?������������������������       �                     �?     @������������������������       �                     �?       @>       m                    �?
�e4���?Q             `@       ?       Z                     �?d�X^_�?I            �\@      *@@       O                    B@H.�!���?!             I@      $@A       N                 `f�D@�LQ�1	�?             7@     @B       C                 ��I*@��S���?
             .@      @������������������������       �                     @        D       E                   �<@z�G�z�?             $@      @������������������������       �                     @      �?F       M                   @>@����X�?             @      @G       L                 �|�?@���Q��?             @       H       I                 �|Y=@�q�q�?             @      @������������������������       �                     �?       J       K                 `fF<@      �?              @      �?������������������������       �                     �?      @������������������������       �                     �?      �?������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        P       Y                 ���[@�����H�?             ;@       Q       X                    �?$�q-�?             :@       R       W                 `f�;@�C��2(�?             6@       S       V                   �K@r�q��?             (@        T       U                 ��:@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@       ������������������������       �                     @        ������������������������       �                     �?        [       l                    �?P�2E��?(            @P@       \       k                   �*@�X�<ݺ?              K@       ]       ^                   �(@$�q-�?            �C@        ������������������������       �        	             ,@        _       `                 �|�<@H%u��?             9@        ������������������������       �                     "@        a       b                 �|�=@     ��?             0@        ������������������������       �                     �?       c       j                   �F@�r����?
             .@       d       i                   @D@z�G�z�?             $@       e       f                    @@�����H�?             "@        ������������������������       �                     @        g       h                   �A@r�q��?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     �?       ������������������������       �                     @       ������������������������       �                     .@       ������������������������       �                     &@       n       o                    :@X�Cc�?             ,@        ������������������������       �                     @        p       q                    5@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        s                          @l���`��?�            �w@       t       �                    �?B�>�;Q�?�            �w@       u       �                    �?C؇eY�?�            �p@        v                        P��@�ucQ?-�?3            @U@        w       ~                 ���@      �?             8@       x       y                 03S@z�G�z�?
             .@        ������������������������       �                     �?       z       {                   �7@d}h���?	             ,@        ������������������������       �                      @        |       }                    �?�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@       ������������������������       �                     "@       �       �                    �?��7��?#            �N@       �       �                 �|Y=@\X��t�?             G@        �       �                    �?     ��?	             0@    p   �       �                   �2@      �?             @    s   ������������������������       �                     �?    f   ������������������������       �                     @        �       �                    �?r�q��?             (@       ������������������������       �                      @        �       �                    ;@      �?             @    n   ������������������������       �                      @        ������������������������       �                      @    o   �       �                    �?�������?             >@    t   ������������������������       �                     @        �       �                 @a'@8����?             7@       �       �                 `�j@�q�q�?             5@   s   �       �                 X��A@�z�G��?             4@   S   �       �                 �;@�����?             3@       �       �                 03@�q�q�?             2@   T   �       �                 ��@�t����?             1@    t   �       �                    �?      �?              @    y   ������������������������       �                     �?    t   ������������������������       �                     �?        �       �                 ���@������?	             .@    ,   ������������������������       �                     �?   y   �       �                    �?����X�?             ,@        ������������������������       �                     @    o   ������������������������       �                     $@       ������������������������       �                     �?    n   ������������������������       �                     �?   m   ������������������������       �                     �?    i   ������������������������       �                     �?       ������������������������       �                      @    e   �       �                    �?z�G�z�?             .@    
   �       �                    &@      �?              @        ������������������������       �                      @   _   ������������������������       �                     @       �       �                 ���&@؇���X�?             @        ������������������������       �                     @    i   �       �                 �|Y=@      �?             @    y   ������������������������       �                     �?        ������������������������       �                     @    n   �       �                   �0@X��Oԣ�?t            @g@    o   ������������������������       �                     @    b   �       �                    �?�8��8��?o            �f@        �       �                 ���@�q�q�?
             .@        ������������������������       �                     �?   t   �       �                 �|�;@����X�?	             ,@       �       �                   �9@���|���?             &@       �       �                    8@�<ݚ�?             "@   l   �       �                   �6@����X�?             @   .   �       �                  �#@r�q��?             @   n   ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @    v   ������������������������       �                     @       �       �                 �?�@�FVQ&�?e            �d@        �       �                 �|Y=@`<)�+�?1            @S@       �       �                   �8@p���?             I@   e   �       �                   �7@ ��WV�?             :@   a   ������������������������       �                     7@        �       �                 `fF@�q�q�?             @    v   ������������������������       �                     �?        ������������������������       �                      @       ������������������������       �                     8@   F   �       �                 �|Y>@�>����?             ;@        �       �                  sW@�t����?
             1@ K@lt ��       �                 ��,@�q�q�?             @    
   ������������������������       �                     @        ������������������������       ��q�q�?             @   ,   ������������������������       �                     &@G   r   ������������������������       �        
             $@       �       �                   �3@`���i��?4             V@    r   �       �                   �1@�θ�?             *@    t   ������������������������       �                      @   c   �       �                 `�8"@���!pc�?             &@       �       �                   �2@և���X�?             @    i   ������������������������       �                     �?    p   ������������������������       ��q�q�?             @    )   ������������������������       �                     @       �       �                   �:@Х-��ٹ?-            �R@    l   ������������������������       �                     <@       �       �                   �;@dP-���?             �G@    t   ������������������������       �                     �?    a   �       �                 @3�@���.�6�?             G@        �       �                   �?@�q�q�?             @    p   ������������������������       �                     �?        ������������������������       �                      @        �       �                 ��) @ �#�Ѵ�?            �E@    t   ������������������������       �                     7@   e   �       �                 �|�>@ףp=
�?             4@       �       �                 pf� @r�q��?
             (@        ������������������������       �                     �?       �       �                    (@�C��2(�?	             &@        �       �                 �|Y=@z�G�z�?             @        �       �                 ���"@      �?              @    t   ������������������������       �                     �?        ������������������������       �                     �?       ������������������������       �                     @       ������������������������       �                     @       ������������������������       �                      @   e   �                          �?������?L             [@   n   �       �                    �?�BE����?)             O@    x   �       �                    �?      �?             $@   i   �       �                    �?X�<ݚ�?             "@       �       �                  S�-@����X�?             @    #   �       �                 03�)@�q�q�?             @    .   ������������������������       �                     �?    t   ������������������������       �                      @    t   ������������������������       �                     @       ������������������������       �                      @        ������������������������       �                     �?   a   �       �                    �?�	j*D�?!             J@   r   �       �                   �3@�P�*�?             ?@        ������������������������       �                     @       �       �                 �|Y=@�q�q�?             ;@        ������������������������       �                     *@   _   �       �                 03�1@X�Cc�?             ,@        �       �                 ���.@ףp=
�?             $@        ������������������������       �                     �?       ������������������������       �                     "@        ������������������������       �                     @    s   �                          �?؇���X�?             5@   a   �                          �?�KM�]�?             3@   r   �                        ��y'@�8��8��?	             (@        �       �                 P�@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                $@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @                                 +@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                 �?*
;&���?#             G@        	                      ��*4@��<b���?             7@        
                        �1@      �?             @        ������������������������       �                      @L \*��                          @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                 @�KM�]�?             3@                                 @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     0@                                 �?���}<S�?             7@       ������������������������       �                     *@                                 @z�G�z�?             $@                              pf�C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                 �?      �?             @        ������������������������       �                     �?                              pf�C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �t�bh�h*h-K ��h/��R�(KMKK��h]�B�       �{@     �p@     �a@     �g@      @      b@      @      K@      @      ?@      @      >@      �?      6@              2@      �?      @      �?                      @      @       @              �?      @      @       @      �?       @                      �?      �?      @              @      �?              @      �?       @              �?      �?              �?      �?                      7@             �V@     �`@     �E@      ;@      4@      3@      3@      1@      &@               @      1@      "@      1@       @      @      @      @      @              @      @                      �?      ,@      @      $@      @      @      @      @      �?       @              �?      �?              �?      �?              �?       @      �?                       @      @              @                      �?       @       @               @       @               @      �?      @              �?      �?              �?      �?             �Z@      7@     @Y@      ,@     �C@      &@      .@       @      @       @      @               @       @              @       @      @       @      @       @      �?      �?              �?      �?      �?                      �?               @               @       @              8@      @      8@       @      4@       @      $@       @      @       @      @                       @      @              $@              @                      �?      O@      @     �I@      @      B@      @      ,@              6@      @      "@              *@      @              �?      *@       @       @       @       @      �?      @              @      �?       @      �?      @                      �?      @              .@              &@              @      "@              @      @       @               @      @              s@     @S@      s@     �R@      l@     �G@     �M@      :@      5@      @      (@      @      �?              &@      @               @      &@      �?              �?      &@              "@              C@      7@      :@      4@      @      *@      �?      @      �?                      @       @      $@               @       @       @       @                       @      7@      @      @              0@      @      ,@      @      ,@      @      *@      @      (@      @      (@      @      �?      �?              �?      �?              &@      @      �?              $@      @              @      $@                      �?      �?              �?                      �?       @              (@      @      @       @               @      @              @      �?      @              @      �?              �?      @             �d@      5@              @     �d@      .@      $@      @              �?      $@      @      @      @      @       @      @       @      @      �?      @                      �?              �?       @                       @      @             `c@      $@     �R@      @     �H@      �?      9@      �?      7@               @      �?              �?       @              8@              9@       @      .@       @      @       @      @              �?       @      &@              $@             @T@      @      $@      @       @               @      @      @      @              �?      @       @      @             �Q@      @      <@             �E@      @              �?     �E@      @       @      �?              �?       @             �D@       @      7@              2@       @      $@       @              �?      $@      �?      @      �?      �?      �?      �?                      �?      @              @               @              T@      <@     �D@      5@      @      @      @      @       @      @       @      �?              �?       @                      @       @              �?              B@      0@      2@      *@              @      2@      "@      *@              @      "@      �?      "@      �?                      "@      @              2@      @      1@       @      &@      �?      @      �?      @                      �?      @              @      �?              �?      @              �?      �?              �?      �?             �C@      @      2@      @      �?      @               @      �?      �?      �?                      �?      1@       @      �?       @      �?                       @      0@              5@       @      *@               @       @      �?       @               @      �?              @               @       @      �?              �?       @               @      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ:9)bhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B�G         �                     @e�L��?�           8�@               Y                     �?x@����?�            �u@               P                   �J@���(�_�?k            �e@y��                          `V�9@�ӭ�a�?Y             b@ ?��  ������������������������       �                     @                                  �7@�:���?T             a@      �?������������������������       �                     3@     �E@       %                   �?@�k��(A�?I            �]@       @	                         x;K@Fx$(�?             I@     "@
                          �<@|��?���?             ;@ ���  ������������������������       �                      @���                            �>@�����?             3@     @                        �|Y=@���Q��?	             .@ ���  ������������������������       �                      @����                            �<@��
ц��?             *@ ���  ������������������������       �                     @���                            @D@���Q��?             $@        ������������������������       �                     @                                  �I@z�G�z�?             @      @������������������������       �                      @       @                           �?�q�q�?             @      @������������������������       �                      @      @������������������������       �                     �?       @������������������������       �                     @               "                    �?��+7��?             7@     �?                           �?�t����?             1@       ������������������������       �                     (@      �?                        `f�N@���Q��?             @      �?������������������������       �                      @     �d@       !                    �?�q�q�?             @      @                          �}S@      �?              @      *@������������������������       �                     �?      "@������������������������       �                     �?        ������������������������       �                     �?      @#       $                    �?�q�q�?             @     �?������������������������       �                     @      @������������������������       �                      @      @&       E                 x5Q@�M���?*             Q@       '       D                 0��M@ҳ�wY;�?             A@       (       1                 ���;@¦	^_�?             ?@      >@)       *                 03k:@8�Z$���?             *@      @������������������������       �                     @       @+       ,                    �?z�G�z�?             $@      @������������������������       �                     �?       @-       .                   �C@�<ݚ�?             "@      �?������������������������       �                     @        /       0                    H@�q�q�?             @     @������������������������       �      �?             @        ������������������������       �                      @        2       5                    �?b�2�tk�?             2@        3       4                 ��A@      �?              @      @������������������������       �                      @        ������������������������       �                     @      �?6       ;                    �?      �?             $@      9@7       :                    �?      �?             @     @8       9                    C@�q�q�?             @      @������������������������       �                      @      &@������������������������       �                     �?        ������������������������       �                     �?        <       =                   �C@      �?             @      0@������������������������       �                     �?       @>       A                    �?���Q��?             @       @?       @                   @A@      �?              @        ������������������������       �                     �?      @������������������������       �                     �?        B       C                 �K@�q�q�?             @      @������������������������       �                      @      �?������������������������       �                     �?       @������������������������       �                     @       @F       G                    �?l��\��?             A@      @������������������������       �        
             0@        H       I                    �?r�q��?	             2@        ������������������������       �                      @        J       O                    �?�z�G��?             $@       K       N                 Ј�U@      �?              @        L       M                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        Q       R                 �U'Q@ܷ��?��?             =@       ������������������������       �                     6@        S       T                    �?և���X�?             @        ������������������������       �                      @        U       V                   �K@z�G�z�?             @        ������������������������       �                      @        W       X                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        Z       _                   �1@և���X�?k            �e@        [       \                    �?�}�+r��?             3@       ������������������������       �                     ,@        ]       ^                    #@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        `       �                    L@����3��?_            �c@       a       |                    �?Fx$(�?Y            �b@        b       {                    :@��ϭ�*�?'             M@       c       d                    �?�����H�?            �F@        ������������������������       �                     @        e       z                    �?,���i�?            �D@       f       s                    �?6YE�t�?            �@@       g       j                   �9@�C��2(�?             6@        h       i                   �3@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        k       l                   �'@�}�+r��?             3@        ������������������������       �                     @        m       r                   �,@�8��8��?             (@       n       o                    B@�����H�?             "@       ������������������������       �                     @        p       q                    D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        t       y                   �E@���!pc�?             &@       u       x                   �;@�����H�?             "@        v       w                   �7@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        
             *@        }       ~                 �|Y=@�nkK�?2             W@        ������������������������       �                     A@               �                   �*@ 	��p�?!             M@       �       �                    �?(N:!���?            �A@        ������������������������       �                     @        �       �                 �|�=@      �?             @@    p   �       �                    @�q�q�?             "@   s   ������������������������       �                     @    f   ������������������������       �                     @        �       �                   @D@�nkK�?             7@       ������������������������       �                     &@        �       �                 `f�)@�8��8��?             (@    n   ������������������������       �                      @        �       �                   �F@ףp=
�?             $@    o   ������������������������       ��q�q�?             @    t   ������������������������       �                     @        ������������������������       �                     7@       ������������������������       �                     @   s   �       �                    @��,?S�?�            �v@    S   �       �                    @$��m��?             :@        ������������������������       �                     &@   T   �       �                    @���Q��?             .@   t   ������������������������       �                     @    y   �       �                    �?      �?              @    t   ������������������������       �                      @        �       �                 ��T?@�q�q�?             @    ,   ������������������������       �                      @   y   ������������������������       �                     @        �       �                    �?�B���?�            u@    o   �       �                   @C@     ��?=             X@       �       �                    �?V�K/��?5            �S@    n   �       �                    �?���B���?             :@   m   �       �                    �?P���Q�?             4@    i   �       �                 ���,@      �?             @       ������������������������       �                     @    e   ������������������������       �                     �?    
   ������������������������       �                     0@        �       �                 `�@1@�q�q�?             @   _   �       �                    �?z�G�z�?             @        ������������������������       �                      @        �       �                 �|Y=@�q�q�?             @    i   ������������������������       �                     �?    y   ������������������������       �                      @        ������������������������       �                     �?    n   �       �                   @A@Fmq��?             �J@   o   �       �                   @1@���Q �?            �H@   b   �       �                    �?)O���?             B@       �       �                   �5@8�A�0��?             6@        �       �                   �3@؇���X�?             @   t   �       �                   !@      �?              @        ������������������������       �                     �?       ������������������������       �                     �?   l   ������������������������       �                     @   .   �       �                 �|�=@��S���?             .@   n   �       �                 ��&@�n_Y�K�?
             *@       �       �                    ;@���!pc�?             &@       �       �                 03�!@և���X�?             @       �       �                   �7@      �?             @        ������������������������       �                      @    v   �       �                 pff@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?       ������������������������       �                     @   e   ������������������������       �                     @   a   ������������������������       �                      @        ������������������������       �                      @    v   �       �                    �?����X�?             ,@       �       �                    �?�θ�?             *@       �       �                 ���)@�q�q�?             "@    F   ������������������������       �                     @        �       �                 �|�;@      �?             @ K@lt �������������������������       �                     �?    
   ������������������������       �                     @        ������������������������       �                     @   ,   ������������������������       �                     �?G   r   ������������������������       �        	             *@       ������������������������       �                     @    r   ������������������������       �                     1@    t   �                          �?P�_��I�?�             n@   c   �       �                    �?      �?�             l@        �       �                 �=/@�<ݚ�?$             K@   i   �       �                   �7@@�0�!��?"            �I@    p   �       �                    �?      �?             @   )   ������������������������       �                      @       ������������������������       �                      @    l   �       �                    �?��0{9�?            �G@        �       �                    �?�X�<ݺ?             2@   t   �       �                 �|Y?@��S�ۿ?             .@   a   �       �                 �|Y;@�����H�?             "@        ������������������������       �                     �?    p   �       �                 ���@      �?              @        ������������������������       �                     @        �       �                 p&�@      �?             @   t   ������������������������       ��q�q�?             @   e   ������������������������       �                     �?       ������������������������       �                     @        ������������������������       �                     @       �       �                  ��@V�a�� �?             =@        ������������������������       �                     @        �       �                    �?���!pc�?             6@   t   �       �                 X��A@����X�?             5@       �       �                   @'@ҳ�wY;�?	             1@       ������������������������       �      �?             0@       ������������������������       �                     �?       ������������������������       �                     @   e   ������������������������       �                     �?   n   ������������������������       �                     @    x   �       �                   �0@��O���?q            @e@    i   �       �                 pf�@      �?             @        ������������������������       �                     �?    #   �       �                    �?���Q��?             @   .   �       �                 pFD!@      �?             @    t   ������������������������       �                      @    t   ������������������������       �                      @       ������������������������       �                     �?        �                         @@@���C"��?l            �d@   a   �                          �? �	.��?V            ``@   r   �                       �!&B@�|K��2�?U             `@       �                       �|�=@�[|x��?S            �_@       �                       �|Y=@@-�_ .�?K            �[@       �                          �?�F��O�?7            @R@   _   �       �                   �:@�U�=���?1            �P@       �       �                 @3�@@9G��?'            �H@       ������������������������       �                     :@       �       �                 0S5 @���}<S�?             7@        �       �                   �2@      �?              @    s   ������������������������       �                     �?   a   �       �                   �3@؇���X�?             @    r   ������������������������       ��q�q�?             @        ������������������������       �                     @       ������������������������       �                     .@                               pf� @@�0�!��?
             1@       ������������������������       �                     "@                             ���)@      �?              @                               �;@      �?             @        ������������������������       �                      @                                �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        	                         5@؇���X�?             @        
                      �Y�@      �?              @        ������������������������       �                     �?sF 5*�� ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     C@                                �?@������?             .@                                �>@      �?              @                              (Se!@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @                              pff@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                 �?؇���X�?             @                             ��I @r�q��?             @       ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                    �@@        ������������������������       �        	             1@        �t�b�(z      h�h*h-K ��h/��R�(KMKK��h]�B�       �{@     �p@     �d@     �f@     �P@     �Z@     �D@     �Y@      @              A@     �Y@              3@      A@      U@      3@      ?@      *@      ,@               @      *@      @      "@      @       @              @      @      @              @      @              @      @      �?       @               @      �?       @                      �?      @              @      1@       @      .@              (@       @      @               @       @      �?      �?      �?              �?      �?              �?              @       @      @                       @      .@     �J@      (@      6@      "@      6@       @      &@              @       @       @              �?       @      @              @       @      @       @       @               @      @      &@       @      @       @                      @      @      @       @       @       @      �?       @                      �?              �?      @      @      �?               @      @      �?      �?              �?      �?              �?       @               @      �?              @              @      ?@              0@      @      .@               @      @      @      �?      @      �?      @              @      �?                      @       @              :@      @      6@              @      @               @      @      �?       @               @      �?              �?       @              Y@     �R@      �?      2@              ,@      �?      @              @      �?             �X@     �L@     @W@     �L@      @     �J@      @      D@              @      @      B@      @      <@       @      4@      �?       @      �?                       @      �?      2@              @      �?      &@      �?       @              @      �?       @      �?                       @              @      @       @      �?       @      �?      @      �?                      @              @       @                       @              *@      V@      @      A@              K@      @      ?@      @      @              <@      @      @      @      @                      @      6@      �?      &@              &@      �?       @              "@      �?       @      �?      @              7@              @             @q@     �U@      "@      1@              &@      "@      @      @               @      @               @       @      @       @                      @     �p@     �Q@      K@      E@     �B@      E@      @      5@      �?      3@      �?      @              @      �?                      0@      @       @      @      �?       @               @      �?              �?       @                      �?      @@      5@      @@      1@      3@      1@      "@      *@      �?      @      �?      �?      �?                      �?              @       @      @       @      @       @      @      @      @      �?      @               @      �?      �?      �?                      �?      @              @                       @               @      $@      @      $@      @      @      @      @              �?      @      �?                      @      @                      �?      *@                      @      1@             �j@      <@     �h@      <@      E@      (@      E@      "@       @       @               @       @              D@      @      1@      �?      ,@      �?       @      �?      �?              @      �?      @              @      �?       @      �?      �?              @              @              7@      @      @              0@      @      .@      @      &@      @      $@      @      �?              @              �?                      @     @c@      0@      @      @      �?               @      @       @       @               @       @                      �?     �b@      *@     �]@      *@      ]@      *@      ]@      $@     @Z@      @     �P@      @     �N@      @     �G@       @      :@              5@       @      @       @              �?      @      �?       @      �?      @              .@              ,@      @      "@              @      @      �?      @               @      �?      �?      �?                      �?      @              @      �?      �?      �?      �?                      �?      @              C@              &@      @      @      @      @       @      @                       @       @      �?       @                      �?      @      �?      @      �?      @      �?       @              �?                      @       @             �@@              1@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�BHzhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMIhuh*h-K ��h/��R�(KMI��h|�B@R         N                    �?�t����?�           8�@     �Y@                           �?�9��L~�?^            �b@      @                        `�@1@�C��2(�?)            �P@      �?                           �?�E��ӭ�?             2@                                  �?�8��8��?             (@       ������������������������       �                     @                                P��+@z�G�z�?             @      @������������������������       �                      @      �?	       
                   �7@�q�q�?             @      @������������������������       �                     �?      @������������������������       �                      @                                   �?�q�q�?             @      @                        �&�)@���Q��?             @        ������������������������       �                     �?                                  �-@      �?             @      �?������������������������       �                      @      &@                        ���,@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?      @������������������������       �                     �?       @                          �H@@��8��?             H@     @������������������������       �                     D@      @                           �?      �?              @       @                           �?      �?             @                               ,w�U@�q�q�?             @      �?������������������������       �                     �?       ������������������������       �                      @      �?������������������������       �                     �?      �?������������������������       �                     @     �d@       -                 pF�#@�t����?5            @U@       @       "                   �5@�#-���?            �A@      *@        !                 �{@      �?              @      "@������������������������       �                     �?        ������������������������       �                     �?      �?#       $                 ���@�FVQ&�?            �@@        ������������������������       �                     ,@      1@%       (                 �|Y=@�KM�]�?             3@      @&       '                   @@      �?             @     @������������������������       �                     @      5@������������������������       �                     �?        )       ,                   @@��S�ۿ?
             .@        *       +                 �|�=@z�G�z�?             @     �?������������������������       �      �?             @      *@������������������������       �                     �?      �?������������������������       �                     $@      @.       I                     @� �	��?             I@     �?/       D                     �?�D����?             E@       0       C                   �H@X�<ݚ�?             B@     @1       2                 �|Y<@���!pc�?             6@        ������������������������       �                     @        3       >                    �?ҳ�wY;�?             1@     <@4       ;                 `f�A@�q�q�?             (@      @5       :                 X�,@@      �?              @     �?6       7                 �ܵ<@���Q��?             @        ������������������������       �                     �?        8       9                 ��2>@      �?             @      @������������������������       �                     @        ������������������������       �                     �?      0@������������������������       �                     @       @<       =                 @�Cq@      �?             @     *@������������������������       �                     @      @������������������������       �                     �?        ?       @                   @H@z�G�z�?             @      �?������������������������       �                     �?      @A       B                    �?      �?             @      @������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     ,@        E       F                 ���@@r�q��?             @     @������������������������       �                     @      �?G       H                    �?      �?              @       @������������������������       �                     �?        ������������������������       �                     �?      �?J       M                    �?      �?              @        K       L                   �3@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        O       �                   �3@�钹H��?^           ��@        P       �                    @��o	��?D             ]@       Q       v                    �?8�$�>�?4            �U@       R       S                    �?
;&����?             G@        ������������������������       �                     @        T       q                    6@�G��l��?             E@       U       n                    �?���Q��?            �A@       V       ]                    �?J�8���?             =@        W       X                   �1@z�G�z�?             @        ������������������������       �                     �?       Y       \                 ��!@      �?             @       Z       [                 P��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ^       a                     @      �?             8@        _       `                   �2@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        b       g                   �1@���y4F�?             3@        c       f                   �0@      �?              @        d       e                 pf�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     @       h       m                 0S5 @���!pc�?             &@        i       j                   �2@      �?             @        ������������������������       �                      @        k       l                 �?�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @       o       p                   �2@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     @        r       s                     �?؇���X�?             @        ������������������������       �                     �?        t       u                   �1@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        w       ~                    �?z�G�z�?             D@        x       y                     @�t����?             1@       ������������������������       �                     $@       z       {                    �?����X�?             @        ������������������������       �                     @        |       }                 `f7@      �?             @       ������������������������       �                      @        ������������������������       �                      @               �                    )@��+7��?             7@       �       �                    �?�KM�]�?             3@       ������������������������       �                     *@       �       �                    �?�q�q�?             @���  �       �                    �?z�G�z�?             @ ���  ������������������������       �                     @ z��  �       �                     �?      �?              @    t   ������������������������       �                     �?    )   ������������������������       �                     �?    e   ������������������������       �                     �?   E   ������������������������       �                     @���  �       �                    �?z�G�z�?             >@ v��  �       �                    @ҳ�wY;�?             1@    e   ������������������������       �                     @��  �       �                    *@��
ц��?             *@   e   �       �                    @�z�G��?             $@        �       �                    @      �?             @    '   ������������������������       �                     �?    x   ������������������������       �                     @����  ������������������������       �                     @   "   ������������������������       �                     @   j   ������������������������       �        	             *@    _   �       �                     @�/e�U��?           �{@ S��  �       �                    �?      �?v             g@��  �       �                    �?*��w\��?\            �b@    s   �       �                    :@=QcG��?            �G@ ���  �       �                   �3@���Q��?             @    p   ������������������������       �                      @ ���  ������������������������       �                     @   e   �       �                   �B@�Ń��̧?             E@��  ������������������������       �                     9@    _   �       �                   @C@�IєX�?             1@    e   ������������������������       �                     �? ���  ������������������������       �        
             0@   t   �       �                    �?��[�8��?B            �Y@    o   ������������������������       �                     �?8��  �       �                     �?�C+����?A            @Y@   m   �       �                    �?���Q �?!            �H@   t   �       �                   �B@�z�G��?             D@   h   �       �                   �A@���Q��?             >@{��  �       �                   �>@�q�q�?             ;@   o   �       �                   @>@և���X�?             5@   x   �       �                 �̌*@�q�q�?             2@    e   ������������������������       �                     @\и�  �       �                 `fF<@և���X�?
             ,@   t   �       �                   @L@�eP*L��?             &@@��  �       �                    H@      �?              @       �       �                 �|�<@      �?             @ ���  ������������������������       �                     �?׸�  �       �                 �|�?@���Q��?             @    n   ������������������������       �                     �?       �       �                   �C@      �?             @ `��  ������������������������       �                     �?�и�  ������������������������       ��q�q�?             @3��  ������������������������       �                      @]   :   ������������������������       �                     @ ���  �       �                 �|Y=@�q�q�?             @    m   ������������������������       �                      @ ��  ������������������������       �                     �?    b   ������������������������       �                     @a��  ������������������������       �                     @ ���  ������������������������       �                     @       ������������������������       �                     $@���  �       �                    =@X�<ݚ�?             "@ ���  ������������������������       �                     �? b��  �       �                 ��<R@      �?              @:��  �       �                   �C@z�G�z�?             @    u   ������������������������       �                      @"   "   �       �                  x#J@�q�q�?             @ U��  ������������������������       �                     �?�T��  �       �                 �K@      �?              @        ������������������������       �                     �?   
   ������������������������       �                     �? Y��  ������������������������       �                     @ Ը�  �       �                    ,@4��?�?              J@���  �       �                 `f�)@�חF�P�?             ?@        ������������������������       �        	             (@�t��  �       �                   �A@�d�����?             3@    r   �       �                 �|Y<@      �?              @ ĸ�  ������������������������       �                      @ |��  �       �                 �|�=@�q�q�?             @ Ǹ�  ������������������������       �                     �?        �       �                    @@���Q��?             @        ������������������������       �                     �?    p   ������������������������       �      �?             @       �       �                   �F@�C��2(�?             &@o��  �       �                   @D@z�G�z�?             @ ��  ������������������������       �                      @ո�  ������������������������       ��q�q�?             @o��  ������������������������       �                     @        ������������������������       �                     5@ ���  �       �                   �M@��R[s�?            �A@:��  �       �                    F@     ��?             @@X��  �       �                    B@�+e�X�?             9@n��  �       �                    �?R���Q�?             4@��  ������������������������       �                     1@���  ������������������������       �                     @    s   �       �                    �?���Q��?             @ i��  ������������������������       �                      @    -   ������������������������       �                     @<���  ������������������������       �                     @   -   ������������������������       �                     @    -   �                          �?�����D�?�            @p@    -   �                          �?�ʻ����?.             Q@ĸ�  �       �                 ��@�~8�e�?$            �I@    c   �       �                    �?@�0�!��?             1@j��  �       �                 ���@ףp=
�?             $@    -   ������������������������       �                     �?    -   ������������������������       �                     "@   -   �       �                 pff@����X�?             @Ǹ�  �       �                 �|�9@      �?             @    m   ������������������������       �                      @       ������������������������       �                      @ ���  ������������������������       �                     @���  �       �                    �?�ʻ����?             A@        ������������������������       �                     @   a   �                         �>@d��0u��?             >@��  �       �                 ��&@l��
I��?             ;@   l   �       �                   �@�r����?
             .@        �       �                 �&B@      �?             @���  �       �                   �7@�q�q�?             @    n   ������������������������       �                     �? ���  ������������������������       �                      @ e��  ������������������������       �                     �?   _   ������������������������       �                     &@   g   �                          4@      �?             (@��  �       �                   �:@      �?              @    r   ������������������������       �                     �? R��  �                           �?؇���X�?             @    r   ������������������������       �                     @    p                           �.@      �?             @        ������������������������       �                     �?       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @                              �|�:@�IєX�?
             1@        ������������������������       �                     �?        ������������������������       �        	             0@        	      D                ���5@     ��?v             h@       
      ?                   �?�L���?r             g@             6                ���"@d#,����?e            �d@@ �*��                          �?@�+9\J�?Z            �b@                              �|Y=@؇���X�?             5@                               ��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                              X�I@�KM�]�?             3@                             ���@�t����?             1@        ������������������������       �                      @                              ��(@�<ݚ�?             "@       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                      @                                �7@����?K            @`@        ������������������������       �                    �A@                              ���@<����?7            �W@        ������������������������       �        	             2@                                @8@�s�c���?.            @S@                              03@      �?             @        ������������������������       �                      @        ������������������������       �                      @               1                @3�@�F��O�?,            @R@       !      "                �|Y=@X�EQ]N�?            �E@        ������������������������       �                     .@        #      0                  �C@�>4և��?             <@       $      %                pf�@�E��ӭ�?             2@        ������������������������       �                     @        &      /                   B@�q�q�?
             (@       '      .                  @@@���|���?	             &@       (      )                  �@���Q��?             $@        ������������������������       �                     @        *      +                �|�>@؇���X�?             @        ������������������������       �                     @        ,      -                �?�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        2      5                �|Y<@(;L]n�?             >@        3      4                  �:@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ;@        7      <                �|�=@d}h���?             ,@       8      9                  �<@�C��2(�?	             &@       ������������������������       �                     @        :      ;                �|Y=@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        =      >                  �A@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        @      C                pf� @P���Q�?             4@        A      B                ��Y@      �?              @       ������������������������       �                     @        ������������������������       �                     �?       ������������������������       �        	             (@       E      H                   �?և���X�?             @        F      G                   �?���Q��?             @        ������������������������       �                      @       ������������������������       �                     @       ������������������������       �                      @       �t�bh�h*h-K ��h/��R�(KMIKK��h]�B�       �z@     �q@     �P@     @U@      @      N@      @      *@      �?      &@              @      �?      @               @      �?       @      �?                       @      @       @      @       @              �?      @      �?       @              �?      �?              �?      �?              �?              �?     �G@              D@      �?      @      �?      @      �?       @      �?                       @              �?              @      N@      9@      @@      @      �?      �?      �?                      �?      ?@       @      ,@              1@       @      @      �?      @                      �?      ,@      �?      @      �?      @      �?      �?              $@              <@      6@      9@      1@      4@      0@      @      0@              @      @      &@      @      @       @      @       @      @      �?              �?      @              @      �?                      @      @      �?      @                      �?      �?      @              �?      �?      @              @      �?              ,@              @      �?      @              �?      �?              �?      �?              @      @      @       @               @      @                      @     `v@     @i@      K@      O@      >@      L@      6@      8@              @      6@      4@      5@      ,@      3@      $@      �?      @              �?      �?      @      �?      �?              �?      �?                       @      2@      @      @       @      @                       @      .@      @      @      �?       @      �?      �?              �?      �?      @               @      @      �?      @               @      �?      �?      �?                      �?      @               @      @       @                      @      �?      @              �?      �?      @      �?                      @       @      @@       @      .@              $@       @      @              @       @       @               @       @              @      1@       @      1@              *@       @      @      �?      @              @      �?      �?      �?                      �?      �?              @              8@      @      &@      @      @              @      @      @      @      �?      @      �?                      @      @                      @      *@              s@     �a@      W@      W@     �T@     �P@      @      F@       @      @       @                      @      �?     �D@              9@      �?      0@      �?                      0@      T@      6@      �?             �S@      6@      @@      1@      <@      (@      2@      (@      2@      "@      (@      "@      (@      @      @               @      @      @      @      @      @      @      @              �?      @       @      �?               @       @              �?       @      �?               @      @               @      �?       @                      �?              @      @                      @      $@              @      @              �?      @      @      @      �?       @               @      �?      �?              �?      �?              �?      �?                      @     �G@      @      :@      @      (@              ,@      @      @      @       @               @      @              �?       @      @      �?              �?      @      $@      �?      @      �?       @               @      �?      @              5@              "@      :@      @      :@      @      3@      @      1@              1@      @              @       @               @      @                      @      @             �j@      H@      C@      >@      6@      =@      @      ,@      �?      "@      �?                      "@       @      @       @       @               @       @                      @      3@      .@              @      3@      &@      3@       @      *@       @       @       @       @      �?              �?       @                      �?      &@              @      @       @      @      �?              �?      @              @      �?      @      �?                      @      @                      @      0@      �?              �?      0@             �e@      2@     @e@      .@     �b@      ,@     �a@      &@      2@      @      �?      �?      �?                      �?      1@       @      .@       @       @              @       @      @       @      �?               @             �^@       @     �A@             �U@       @      2@             @Q@       @       @       @               @       @             �P@      @      C@      @      .@              7@      @      *@      @      @              @      @      @      @      @      @              @      @      �?      @               @      �?      �?              �?      �?      �?                      �?      $@              =@      �?       @      �?       @                      �?      ;@              &@      @      $@      �?      @              @      �?              �?      @              �?       @               @      �?              3@      �?      @      �?      @                      �?      (@              @      @       @      @       @                      @       @        �t�bubhhubehhub.